netcdf temp_year { 
dimensions:
    time_temp_year = 8761;
    temp_year = 8761;

variables:

    double temp_year(time_temp_year) ;
        temp_year:interpolation = "discrete" ;

    double time_temp_year(time_temp_year) ;
        time_temp_year:extrapolation = "periodic" ;
        time_temp_year:add_offset = 0.f;
//global attributes:
:float_ex=1.1f;
:TRY=2010;
:Region=12;
data:

     time_temp_year=
        0.0, 3600.0, 7200.0, 10800.0, 14400.0, 18000.0, 21600.0, 25200.0, 28800.0, 32400.0, 36000.0, 39600.0, 43200.0, 46800.0, 50400.0, 54000.0, 57600.0, 61200.0, 64800.0, 68400.0, 72000.0, 75600.0, 79200.0, 82800.0, 86400.0, 90000.0, 93600.0, 97200.0, 100800.0, 104400.0, 108000.0, 111600.0, 115200.0, 118800.0, 122400.0, 126000.0, 129600.0, 133200.0, 136800.0, 140400.0, 144000.0, 147600.0, 151200.0, 154800.0, 158400.0, 162000.0, 165600.0, 169200.0, 172800.0, 176400.0, 180000.0, 183600.0, 187200.0, 190800.0, 194400.0, 198000.0, 201600.0, 205200.0, 208800.0, 212400.0, 216000.0, 219600.0, 223200.0, 226800.0, 230400.0, 234000.0, 237600.0, 241200.0, 244800.0, 248400.0, 252000.0, 255600.0, 259200.0, 262800.0, 266400.0, 270000.0, 273600.0, 277200.0, 280800.0, 284400.0, 288000.0, 291600.0, 295200.0, 298800.0, 302400.0, 306000.0, 309600.0, 313200.0, 316800.0, 320400.0, 324000.0, 327600.0, 331200.0, 334800.0, 338400.0, 342000.0, 345600.0, 349200.0, 352800.0, 356400.0, 360000.0, 363600.0, 367200.0, 370800.0, 374400.0, 378000.0, 381600.0, 385200.0, 388800.0, 392400.0, 396000.0, 399600.0, 403200.0, 406800.0, 410400.0, 414000.0, 417600.0, 421200.0, 424800.0, 428400.0, 432000.0, 435600.0, 439200.0, 442800.0, 446400.0, 450000.0, 453600.0, 457200.0, 460800.0, 464400.0, 468000.0, 471600.0, 475200.0, 478800.0, 482400.0, 486000.0, 489600.0, 493200.0, 496800.0, 500400.0, 504000.0, 507600.0, 511200.0, 514800.0, 518400.0, 522000.0, 525600.0, 529200.0, 532800.0, 536400.0, 540000.0, 543600.0, 547200.0, 550800.0, 554400.0, 558000.0, 561600.0, 565200.0, 568800.0, 572400.0, 576000.0, 579600.0, 583200.0, 586800.0, 590400.0, 594000.0, 597600.0, 601200.0, 604800.0, 608400.0, 612000.0, 615600.0, 619200.0, 622800.0, 626400.0, 630000.0, 633600.0, 637200.0, 640800.0, 644400.0, 648000.0, 651600.0, 655200.0, 658800.0, 662400.0, 666000.0, 669600.0, 673200.0, 676800.0, 680400.0, 684000.0, 687600.0, 691200.0, 694800.0, 698400.0, 702000.0, 705600.0, 709200.0, 712800.0, 716400.0, 720000.0, 723600.0, 727200.0, 730800.0, 734400.0, 738000.0, 741600.0, 745200.0, 748800.0, 752400.0, 756000.0, 759600.0, 763200.0, 766800.0, 770400.0, 774000.0, 777600.0, 781200.0, 784800.0, 788400.0, 792000.0, 795600.0, 799200.0, 802800.0, 806400.0, 810000.0, 813600.0, 817200.0, 820800.0, 824400.0, 828000.0, 831600.0, 835200.0, 838800.0, 842400.0, 846000.0, 849600.0, 853200.0, 856800.0, 860400.0, 864000.0, 867600.0, 871200.0, 874800.0, 878400.0, 882000.0, 885600.0, 889200.0, 892800.0, 896400.0, 900000.0, 903600.0, 907200.0, 910800.0, 914400.0, 918000.0, 921600.0, 925200.0, 928800.0, 932400.0, 936000.0, 939600.0, 943200.0, 946800.0, 950400.0, 954000.0, 957600.0, 961200.0, 964800.0, 968400.0, 972000.0, 975600.0, 979200.0, 982800.0, 986400.0, 990000.0, 993600.0, 997200.0, 1000800.0, 1004400.0, 1008000.0, 1011600.0, 1015200.0, 1018800.0, 1022400.0, 1026000.0, 1029600.0, 1033200.0, 1036800.0, 1040400.0, 1044000.0, 1047600.0, 1051200.0, 1054800.0, 1058400.0, 1062000.0, 1065600.0, 1069200.0, 1072800.0, 1076400.0, 1080000.0, 1083600.0, 1087200.0, 1090800.0, 1094400.0, 1098000.0, 1101600.0, 1105200.0, 1108800.0, 1112400.0, 1116000.0, 1119600.0, 1123200.0, 1126800.0, 1130400.0, 1134000.0, 1137600.0, 1141200.0, 1144800.0, 1148400.0, 1152000.0, 1155600.0, 1159200.0, 1162800.0, 1166400.0, 1170000.0, 1173600.0, 1177200.0, 1180800.0, 1184400.0, 1188000.0, 1191600.0, 1195200.0, 1198800.0, 1202400.0, 1206000.0, 1209600.0, 1213200.0, 1216800.0, 1220400.0, 1224000.0, 1227600.0, 1231200.0, 1234800.0, 1238400.0, 1242000.0, 1245600.0, 1249200.0, 1252800.0, 1256400.0, 1260000.0, 1263600.0, 1267200.0, 1270800.0, 1274400.0, 1278000.0, 1281600.0, 1285200.0, 1288800.0, 1292400.0, 1296000.0, 1299600.0, 1303200.0, 1306800.0, 1310400.0, 1314000.0, 1317600.0, 1321200.0, 1324800.0, 1328400.0, 1332000.0, 1335600.0, 1339200.0, 1342800.0, 1346400.0, 1350000.0, 1353600.0, 1357200.0, 1360800.0, 1364400.0, 1368000.0, 1371600.0, 1375200.0, 1378800.0, 1382400.0, 1386000.0, 1389600.0, 1393200.0, 1396800.0, 1400400.0, 1404000.0, 1407600.0, 1411200.0, 1414800.0, 1418400.0, 1422000.0, 1425600.0, 1429200.0, 1432800.0, 1436400.0, 1440000.0, 1443600.0, 1447200.0, 1450800.0, 1454400.0, 1458000.0, 1461600.0, 1465200.0, 1468800.0, 1472400.0, 1476000.0, 1479600.0, 1483200.0, 1486800.0, 1490400.0, 1494000.0, 1497600.0, 1501200.0, 1504800.0, 1508400.0, 1512000.0, 1515600.0, 1519200.0, 1522800.0, 1526400.0, 1530000.0, 1533600.0, 1537200.0, 1540800.0, 1544400.0, 1548000.0, 1551600.0, 1555200.0, 1558800.0, 1562400.0, 1566000.0, 1569600.0, 1573200.0, 1576800.0, 1580400.0, 1584000.0, 1587600.0, 1591200.0, 1594800.0, 1598400.0, 1602000.0, 1605600.0, 1609200.0, 1612800.0, 1616400.0, 1620000.0, 1623600.0, 1627200.0, 1630800.0, 1634400.0, 1638000.0, 1641600.0, 1645200.0, 1648800.0, 1652400.0, 1656000.0, 1659600.0, 1663200.0, 1666800.0, 1670400.0, 1674000.0, 1677600.0, 1681200.0, 1684800.0, 1688400.0, 1692000.0, 1695600.0, 1699200.0, 1702800.0, 1706400.0, 1710000.0, 1713600.0, 1717200.0, 1720800.0, 1724400.0, 1728000.0, 1731600.0, 1735200.0, 1738800.0, 1742400.0, 1746000.0, 1749600.0, 1753200.0, 1756800.0, 1760400.0, 1764000.0, 1767600.0, 1771200.0, 1774800.0, 1778400.0, 1782000.0, 1785600.0, 1789200.0, 1792800.0, 1796400.0, 1800000.0, 1803600.0, 1807200.0, 1810800.0, 1814400.0, 1818000.0, 1821600.0, 1825200.0, 1828800.0, 1832400.0, 1836000.0, 1839600.0, 1843200.0, 1846800.0, 1850400.0, 1854000.0, 1857600.0, 1861200.0, 1864800.0, 1868400.0, 1872000.0, 1875600.0, 1879200.0, 1882800.0, 1886400.0, 1890000.0, 1893600.0, 1897200.0, 1900800.0, 1904400.0, 1908000.0, 1911600.0, 1915200.0, 1918800.0, 1922400.0, 1926000.0, 1929600.0, 1933200.0, 1936800.0, 1940400.0, 1944000.0, 1947600.0, 1951200.0, 1954800.0, 1958400.0, 1962000.0, 1965600.0, 1969200.0, 1972800.0, 1976400.0, 1980000.0, 1983600.0, 1987200.0, 1990800.0, 1994400.0, 1998000.0, 2001600.0, 2005200.0, 2008800.0, 2012400.0, 2016000.0, 2019600.0, 2023200.0, 2026800.0, 2030400.0, 2034000.0, 2037600.0, 2041200.0, 2044800.0, 2048400.0, 2052000.0, 2055600.0, 2059200.0, 2062800.0, 2066400.0, 2070000.0, 2073600.0, 2077200.0, 2080800.0, 2084400.0, 2088000.0, 2091600.0, 2095200.0, 2098800.0, 2102400.0, 2106000.0, 2109600.0, 2113200.0, 2116800.0, 2120400.0, 2124000.0, 2127600.0, 2131200.0, 2134800.0, 2138400.0, 2142000.0, 2145600.0, 2149200.0, 2152800.0, 2156400.0, 2160000.0, 2163600.0, 2167200.0, 2170800.0, 2174400.0, 2178000.0, 2181600.0, 2185200.0, 2188800.0, 2192400.0, 2196000.0, 2199600.0, 2203200.0, 2206800.0, 2210400.0, 2214000.0, 2217600.0, 2221200.0, 2224800.0, 2228400.0, 2232000.0, 2235600.0, 2239200.0, 2242800.0, 2246400.0, 2250000.0, 2253600.0, 2257200.0, 2260800.0, 2264400.0, 2268000.0, 2271600.0, 2275200.0, 2278800.0, 2282400.0, 2286000.0, 2289600.0, 2293200.0, 2296800.0, 2300400.0, 2304000.0, 2307600.0, 2311200.0, 2314800.0, 2318400.0, 2322000.0, 2325600.0, 2329200.0, 2332800.0, 2336400.0, 2340000.0, 2343600.0, 2347200.0, 2350800.0, 2354400.0, 2358000.0, 2361600.0, 2365200.0, 2368800.0, 2372400.0, 2376000.0, 2379600.0, 2383200.0, 2386800.0, 2390400.0, 2394000.0, 2397600.0, 2401200.0, 2404800.0, 2408400.0, 2412000.0, 2415600.0, 2419200.0, 2422800.0, 2426400.0, 2430000.0, 2433600.0, 2437200.0, 2440800.0, 2444400.0, 2448000.0, 2451600.0, 2455200.0, 2458800.0, 2462400.0, 2466000.0, 2469600.0, 2473200.0, 2476800.0, 2480400.0, 2484000.0, 2487600.0, 2491200.0, 2494800.0, 2498400.0, 2502000.0, 2505600.0, 2509200.0, 2512800.0, 2516400.0, 2520000.0, 2523600.0, 2527200.0, 2530800.0, 2534400.0, 2538000.0, 2541600.0, 2545200.0, 2548800.0, 2552400.0, 2556000.0, 2559600.0, 2563200.0, 2566800.0, 2570400.0, 2574000.0, 2577600.0, 2581200.0, 2584800.0, 2588400.0, 2592000.0, 2595600.0, 2599200.0, 2602800.0, 2606400.0, 2610000.0, 2613600.0, 2617200.0, 2620800.0, 2624400.0, 2628000.0, 2631600.0, 2635200.0, 2638800.0, 2642400.0, 2646000.0, 2649600.0, 2653200.0, 2656800.0, 2660400.0, 2664000.0, 2667600.0, 2671200.0, 2674800.0, 2678400.0, 2682000.0, 2685600.0, 2689200.0, 2692800.0, 2696400.0, 2700000.0, 2703600.0, 2707200.0, 2710800.0, 2714400.0, 2718000.0, 2721600.0, 2725200.0, 2728800.0, 2732400.0, 2736000.0, 2739600.0, 2743200.0, 2746800.0, 2750400.0, 2754000.0, 2757600.0, 2761200.0, 2764800.0, 2768400.0, 2772000.0, 2775600.0, 2779200.0, 2782800.0, 2786400.0, 2790000.0, 2793600.0, 2797200.0, 2800800.0, 2804400.0, 2808000.0, 2811600.0, 2815200.0, 2818800.0, 2822400.0, 2826000.0, 2829600.0, 2833200.0, 2836800.0, 2840400.0, 2844000.0, 2847600.0, 2851200.0, 2854800.0, 2858400.0, 2862000.0, 2865600.0, 2869200.0, 2872800.0, 2876400.0, 2880000.0, 2883600.0, 2887200.0, 2890800.0, 2894400.0, 2898000.0, 2901600.0, 2905200.0, 2908800.0, 2912400.0, 2916000.0, 2919600.0, 2923200.0, 2926800.0, 2930400.0, 2934000.0, 2937600.0, 2941200.0, 2944800.0, 2948400.0, 2952000.0, 2955600.0, 2959200.0, 2962800.0, 2966400.0, 2970000.0, 2973600.0, 2977200.0, 2980800.0, 2984400.0, 2988000.0, 2991600.0, 2995200.0, 2998800.0, 3002400.0, 3006000.0, 3009600.0, 3013200.0, 3016800.0, 3020400.0, 3024000.0, 3027600.0, 3031200.0, 3034800.0, 3038400.0, 3042000.0, 3045600.0, 3049200.0, 3052800.0, 3056400.0, 3060000.0, 3063600.0, 3067200.0, 3070800.0, 3074400.0, 3078000.0, 3081600.0, 3085200.0, 3088800.0, 3092400.0, 3096000.0, 3099600.0, 3103200.0, 3106800.0, 3110400.0, 3114000.0, 3117600.0, 3121200.0, 3124800.0, 3128400.0, 3132000.0, 3135600.0, 3139200.0, 3142800.0, 3146400.0, 3150000.0, 3153600.0, 3157200.0, 3160800.0, 3164400.0, 3168000.0, 3171600.0, 3175200.0, 3178800.0, 3182400.0, 3186000.0, 3189600.0, 3193200.0, 3196800.0, 3200400.0, 3204000.0, 3207600.0, 3211200.0, 3214800.0, 3218400.0, 3222000.0, 3225600.0, 3229200.0, 3232800.0, 3236400.0, 3240000.0, 3243600.0, 3247200.0, 3250800.0, 3254400.0, 3258000.0, 3261600.0, 3265200.0, 3268800.0, 3272400.0, 3276000.0, 3279600.0, 3283200.0, 3286800.0, 3290400.0, 3294000.0, 3297600.0, 3301200.0, 3304800.0, 3308400.0, 3312000.0, 3315600.0, 3319200.0, 3322800.0, 3326400.0, 3330000.0, 3333600.0, 3337200.0, 3340800.0, 3344400.0, 3348000.0, 3351600.0, 3355200.0, 3358800.0, 3362400.0, 3366000.0, 3369600.0, 3373200.0, 3376800.0, 3380400.0, 3384000.0, 3387600.0, 3391200.0, 3394800.0, 3398400.0, 3402000.0, 3405600.0, 3409200.0, 3412800.0, 3416400.0, 3420000.0, 3423600.0, 3427200.0, 3430800.0, 3434400.0, 3438000.0, 3441600.0, 3445200.0, 3448800.0, 3452400.0, 3456000.0, 3459600.0, 3463200.0, 3466800.0, 3470400.0, 3474000.0, 3477600.0, 3481200.0, 3484800.0, 3488400.0, 3492000.0, 3495600.0, 3499200.0, 3502800.0, 3506400.0, 3510000.0, 3513600.0, 3517200.0, 3520800.0, 3524400.0, 3528000.0, 3531600.0, 3535200.0, 3538800.0, 3542400.0, 3546000.0, 3549600.0, 3553200.0, 3556800.0, 3560400.0, 3564000.0, 3567600.0, 3571200.0, 3574800.0, 3578400.0, 3582000.0, 3585600.0, 3589200.0, 3592800.0, 3596400.0, 3600000.0, 3603600.0, 3607200.0, 3610800.0, 3614400.0, 3618000.0, 3621600.0, 3625200.0, 3628800.0, 3632400.0, 3636000.0, 3639600.0, 3643200.0, 3646800.0, 3650400.0, 3654000.0, 3657600.0, 3661200.0, 3664800.0, 3668400.0, 3672000.0, 3675600.0, 3679200.0, 3682800.0, 3686400.0, 3690000.0, 3693600.0, 3697200.0, 3700800.0, 3704400.0, 3708000.0, 3711600.0, 3715200.0, 3718800.0, 3722400.0, 3726000.0, 3729600.0, 3733200.0, 3736800.0, 3740400.0, 3744000.0, 3747600.0, 3751200.0, 3754800.0, 3758400.0, 3762000.0, 3765600.0, 3769200.0, 3772800.0, 3776400.0, 3780000.0, 3783600.0, 3787200.0, 3790800.0, 3794400.0, 3798000.0, 3801600.0, 3805200.0, 3808800.0, 3812400.0, 3816000.0, 3819600.0, 3823200.0, 3826800.0, 3830400.0, 3834000.0, 3837600.0, 3841200.0, 3844800.0, 3848400.0, 3852000.0, 3855600.0, 3859200.0, 3862800.0, 3866400.0, 3870000.0, 3873600.0, 3877200.0, 3880800.0, 3884400.0, 3888000.0, 3891600.0, 3895200.0, 3898800.0, 3902400.0, 3906000.0, 3909600.0, 3913200.0, 3916800.0, 3920400.0, 3924000.0, 3927600.0, 3931200.0, 3934800.0, 3938400.0, 3942000.0, 3945600.0, 3949200.0, 3952800.0, 3956400.0, 3960000.0, 3963600.0, 3967200.0, 3970800.0, 3974400.0, 3978000.0, 3981600.0, 3985200.0, 3988800.0, 3992400.0, 3996000.0, 3999600.0, 4003200.0, 4006800.0, 4010400.0, 4014000.0, 4017600.0, 4021200.0, 4024800.0, 4028400.0, 4032000.0, 4035600.0, 4039200.0, 4042800.0, 4046400.0, 4050000.0, 4053600.0, 4057200.0, 4060800.0, 4064400.0, 4068000.0, 4071600.0, 4075200.0, 4078800.0, 4082400.0, 4086000.0, 4089600.0, 4093200.0, 4096800.0, 4100400.0, 4104000.0, 4107600.0, 4111200.0, 4114800.0, 4118400.0, 4122000.0, 4125600.0, 4129200.0, 4132800.0, 4136400.0, 4140000.0, 4143600.0, 4147200.0, 4150800.0, 4154400.0, 4158000.0, 4161600.0, 4165200.0, 4168800.0, 4172400.0, 4176000.0, 4179600.0, 4183200.0, 4186800.0, 4190400.0, 4194000.0, 4197600.0, 4201200.0, 4204800.0, 4208400.0, 4212000.0, 4215600.0, 4219200.0, 4222800.0, 4226400.0, 4230000.0, 4233600.0, 4237200.0, 4240800.0, 4244400.0, 4248000.0, 4251600.0, 4255200.0, 4258800.0, 4262400.0, 4266000.0, 4269600.0, 4273200.0, 4276800.0, 4280400.0, 4284000.0, 4287600.0, 4291200.0, 4294800.0, 4298400.0, 4302000.0, 4305600.0, 4309200.0, 4312800.0, 4316400.0, 4320000.0, 4323600.0, 4327200.0, 4330800.0, 4334400.0, 4338000.0, 4341600.0, 4345200.0, 4348800.0, 4352400.0, 4356000.0, 4359600.0, 4363200.0, 4366800.0, 4370400.0, 4374000.0, 4377600.0, 4381200.0, 4384800.0, 4388400.0, 4392000.0, 4395600.0, 4399200.0, 4402800.0, 4406400.0, 4410000.0, 4413600.0, 4417200.0, 4420800.0, 4424400.0, 4428000.0, 4431600.0, 4435200.0, 4438800.0, 4442400.0, 4446000.0, 4449600.0, 4453200.0, 4456800.0, 4460400.0, 4464000.0, 4467600.0, 4471200.0, 4474800.0, 4478400.0, 4482000.0, 4485600.0, 4489200.0, 4492800.0, 4496400.0, 4500000.0, 4503600.0, 4507200.0, 4510800.0, 4514400.0, 4518000.0, 4521600.0, 4525200.0, 4528800.0, 4532400.0, 4536000.0, 4539600.0, 4543200.0, 4546800.0, 4550400.0, 4554000.0, 4557600.0, 4561200.0, 4564800.0, 4568400.0, 4572000.0, 4575600.0, 4579200.0, 4582800.0, 4586400.0, 4590000.0, 4593600.0, 4597200.0, 4600800.0, 4604400.0, 4608000.0, 4611600.0, 4615200.0, 4618800.0, 4622400.0, 4626000.0, 4629600.0, 4633200.0, 4636800.0, 4640400.0, 4644000.0, 4647600.0, 4651200.0, 4654800.0, 4658400.0, 4662000.0, 4665600.0, 4669200.0, 4672800.0, 4676400.0, 4680000.0, 4683600.0, 4687200.0, 4690800.0, 4694400.0, 4698000.0, 4701600.0, 4705200.0, 4708800.0, 4712400.0, 4716000.0, 4719600.0, 4723200.0, 4726800.0, 4730400.0, 4734000.0, 4737600.0, 4741200.0, 4744800.0, 4748400.0, 4752000.0, 4755600.0, 4759200.0, 4762800.0, 4766400.0, 4770000.0, 4773600.0, 4777200.0, 4780800.0, 4784400.0, 4788000.0, 4791600.0, 4795200.0, 4798800.0, 4802400.0, 4806000.0, 4809600.0, 4813200.0, 4816800.0, 4820400.0, 4824000.0, 4827600.0, 4831200.0, 4834800.0, 4838400.0, 4842000.0, 4845600.0, 4849200.0, 4852800.0, 4856400.0, 4860000.0, 4863600.0, 4867200.0, 4870800.0, 4874400.0, 4878000.0, 4881600.0, 4885200.0, 4888800.0, 4892400.0, 4896000.0, 4899600.0, 4903200.0, 4906800.0, 4910400.0, 4914000.0, 4917600.0, 4921200.0, 4924800.0, 4928400.0, 4932000.0, 4935600.0, 4939200.0, 4942800.0, 4946400.0, 4950000.0, 4953600.0, 4957200.0, 4960800.0, 4964400.0, 4968000.0, 4971600.0, 4975200.0, 4978800.0, 4982400.0, 4986000.0, 4989600.0, 4993200.0, 4996800.0, 5000400.0, 5004000.0, 5007600.0, 5011200.0, 5014800.0, 5018400.0, 5022000.0, 5025600.0, 5029200.0, 5032800.0, 5036400.0, 5040000.0, 5043600.0, 5047200.0, 5050800.0, 5054400.0, 5058000.0, 5061600.0, 5065200.0, 5068800.0, 5072400.0, 5076000.0, 5079600.0, 5083200.0, 5086800.0, 5090400.0, 5094000.0, 5097600.0, 5101200.0, 5104800.0, 5108400.0, 5112000.0, 5115600.0, 5119200.0, 5122800.0, 5126400.0, 5130000.0, 5133600.0, 5137200.0, 5140800.0, 5144400.0, 5148000.0, 5151600.0, 5155200.0, 5158800.0, 5162400.0, 5166000.0, 5169600.0, 5173200.0, 5176800.0, 5180400.0, 5184000.0, 5187600.0, 5191200.0, 5194800.0, 5198400.0, 5202000.0, 5205600.0, 5209200.0, 5212800.0, 5216400.0, 5220000.0, 5223600.0, 5227200.0, 5230800.0, 5234400.0, 5238000.0, 5241600.0, 5245200.0, 5248800.0, 5252400.0, 5256000.0, 5259600.0, 5263200.0, 5266800.0, 5270400.0, 5274000.0, 5277600.0, 5281200.0, 5284800.0, 5288400.0, 5292000.0, 5295600.0, 5299200.0, 5302800.0, 5306400.0, 5310000.0, 5313600.0, 5317200.0, 5320800.0, 5324400.0, 5328000.0, 5331600.0, 5335200.0, 5338800.0, 5342400.0, 5346000.0, 5349600.0, 5353200.0, 5356800.0, 5360400.0, 5364000.0, 5367600.0, 5371200.0, 5374800.0, 5378400.0, 5382000.0, 5385600.0, 5389200.0, 5392800.0, 5396400.0, 5400000.0, 5403600.0, 5407200.0, 5410800.0, 5414400.0, 5418000.0, 5421600.0, 5425200.0, 5428800.0, 5432400.0, 5436000.0, 5439600.0, 5443200.0, 5446800.0, 5450400.0, 5454000.0, 5457600.0, 5461200.0, 5464800.0, 5468400.0, 5472000.0, 5475600.0, 5479200.0, 5482800.0, 5486400.0, 5490000.0, 5493600.0, 5497200.0, 5500800.0, 5504400.0, 5508000.0, 5511600.0, 5515200.0, 5518800.0, 5522400.0, 5526000.0, 5529600.0, 5533200.0, 5536800.0, 5540400.0, 5544000.0, 5547600.0, 5551200.0, 5554800.0, 5558400.0, 5562000.0, 5565600.0, 5569200.0, 5572800.0, 5576400.0, 5580000.0, 5583600.0, 5587200.0, 5590800.0, 5594400.0, 5598000.0, 5601600.0, 5605200.0, 5608800.0, 5612400.0, 5616000.0, 5619600.0, 5623200.0, 5626800.0, 5630400.0, 5634000.0, 5637600.0, 5641200.0, 5644800.0, 5648400.0, 5652000.0, 5655600.0, 5659200.0, 5662800.0, 5666400.0, 5670000.0, 5673600.0, 5677200.0, 5680800.0, 5684400.0, 5688000.0, 5691600.0, 5695200.0, 5698800.0, 5702400.0, 5706000.0, 5709600.0, 5713200.0, 5716800.0, 5720400.0, 5724000.0, 5727600.0, 5731200.0, 5734800.0, 5738400.0, 5742000.0, 5745600.0, 5749200.0, 5752800.0, 5756400.0, 5760000.0, 5763600.0, 5767200.0, 5770800.0, 5774400.0, 5778000.0, 5781600.0, 5785200.0, 5788800.0, 5792400.0, 5796000.0, 5799600.0, 5803200.0, 5806800.0, 5810400.0, 5814000.0, 5817600.0, 5821200.0, 5824800.0, 5828400.0, 5832000.0, 5835600.0, 5839200.0, 5842800.0, 5846400.0, 5850000.0, 5853600.0, 5857200.0, 5860800.0, 5864400.0, 5868000.0, 5871600.0, 5875200.0, 5878800.0, 5882400.0, 5886000.0, 5889600.0, 5893200.0, 5896800.0, 5900400.0, 5904000.0, 5907600.0, 5911200.0, 5914800.0, 5918400.0, 5922000.0, 5925600.0, 5929200.0, 5932800.0, 5936400.0, 5940000.0, 5943600.0, 5947200.0, 5950800.0, 5954400.0, 5958000.0, 5961600.0, 5965200.0, 5968800.0, 5972400.0, 5976000.0, 5979600.0, 5983200.0, 5986800.0, 5990400.0, 5994000.0, 5997600.0, 6001200.0, 6004800.0, 6008400.0, 6012000.0, 6015600.0, 6019200.0, 6022800.0, 6026400.0, 6030000.0, 6033600.0, 6037200.0, 6040800.0, 6044400.0, 6048000.0, 6051600.0, 6055200.0, 6058800.0, 6062400.0, 6066000.0, 6069600.0, 6073200.0, 6076800.0, 6080400.0, 6084000.0, 6087600.0, 6091200.0, 6094800.0, 6098400.0, 6102000.0, 6105600.0, 6109200.0, 6112800.0, 6116400.0, 6120000.0, 6123600.0, 6127200.0, 6130800.0, 6134400.0, 6138000.0, 6141600.0, 6145200.0, 6148800.0, 6152400.0, 6156000.0, 6159600.0, 6163200.0, 6166800.0, 6170400.0, 6174000.0, 6177600.0, 6181200.0, 6184800.0, 6188400.0, 6192000.0, 6195600.0, 6199200.0, 6202800.0, 6206400.0, 6210000.0, 6213600.0, 6217200.0, 6220800.0, 6224400.0, 6228000.0, 6231600.0, 6235200.0, 6238800.0, 6242400.0, 6246000.0, 6249600.0, 6253200.0, 6256800.0, 6260400.0, 6264000.0, 6267600.0, 6271200.0, 6274800.0, 6278400.0, 6282000.0, 6285600.0, 6289200.0, 6292800.0, 6296400.0, 6300000.0, 6303600.0, 6307200.0, 6310800.0, 6314400.0, 6318000.0, 6321600.0, 6325200.0, 6328800.0, 6332400.0, 6336000.0, 6339600.0, 6343200.0, 6346800.0, 6350400.0, 6354000.0, 6357600.0, 6361200.0, 6364800.0, 6368400.0, 6372000.0, 6375600.0, 6379200.0, 6382800.0, 6386400.0, 6390000.0, 6393600.0, 6397200.0, 6400800.0, 6404400.0, 6408000.0, 6411600.0, 6415200.0, 6418800.0, 6422400.0, 6426000.0, 6429600.0, 6433200.0, 6436800.0, 6440400.0, 6444000.0, 6447600.0, 6451200.0, 6454800.0, 6458400.0, 6462000.0, 6465600.0, 6469200.0, 6472800.0, 6476400.0, 6480000.0, 6483600.0, 6487200.0, 6490800.0, 6494400.0, 6498000.0, 6501600.0, 6505200.0, 6508800.0, 6512400.0, 6516000.0, 6519600.0, 6523200.0, 6526800.0, 6530400.0, 6534000.0, 6537600.0, 6541200.0, 6544800.0, 6548400.0, 6552000.0, 6555600.0, 6559200.0, 6562800.0, 6566400.0, 6570000.0, 6573600.0, 6577200.0, 6580800.0, 6584400.0, 6588000.0, 6591600.0, 6595200.0, 6598800.0, 6602400.0, 6606000.0, 6609600.0, 6613200.0, 6616800.0, 6620400.0, 6624000.0, 6627600.0, 6631200.0, 6634800.0, 6638400.0, 6642000.0, 6645600.0, 6649200.0, 6652800.0, 6656400.0, 6660000.0, 6663600.0, 6667200.0, 6670800.0, 6674400.0, 6678000.0, 6681600.0, 6685200.0, 6688800.0, 6692400.0, 6696000.0, 6699600.0, 6703200.0, 6706800.0, 6710400.0, 6714000.0, 6717600.0, 6721200.0, 6724800.0, 6728400.0, 6732000.0, 6735600.0, 6739200.0, 6742800.0, 6746400.0, 6750000.0, 6753600.0, 6757200.0, 6760800.0, 6764400.0, 6768000.0, 6771600.0, 6775200.0, 6778800.0, 6782400.0, 6786000.0, 6789600.0, 6793200.0, 6796800.0, 6800400.0, 6804000.0, 6807600.0, 6811200.0, 6814800.0, 6818400.0, 6822000.0, 6825600.0, 6829200.0, 6832800.0, 6836400.0, 6840000.0, 6843600.0, 6847200.0, 6850800.0, 6854400.0, 6858000.0, 6861600.0, 6865200.0, 6868800.0, 6872400.0, 6876000.0, 6879600.0, 6883200.0, 6886800.0, 6890400.0, 6894000.0, 6897600.0, 6901200.0, 6904800.0, 6908400.0, 6912000.0, 6915600.0, 6919200.0, 6922800.0, 6926400.0, 6930000.0, 6933600.0, 6937200.0, 6940800.0, 6944400.0, 6948000.0, 6951600.0, 6955200.0, 6958800.0, 6962400.0, 6966000.0, 6969600.0, 6973200.0, 6976800.0, 6980400.0, 6984000.0, 6987600.0, 6991200.0, 6994800.0, 6998400.0, 7002000.0, 7005600.0, 7009200.0, 7012800.0, 7016400.0, 7020000.0, 7023600.0, 7027200.0, 7030800.0, 7034400.0, 7038000.0, 7041600.0, 7045200.0, 7048800.0, 7052400.0, 7056000.0, 7059600.0, 7063200.0, 7066800.0, 7070400.0, 7074000.0, 7077600.0, 7081200.0, 7084800.0, 7088400.0, 7092000.0, 7095600.0, 7099200.0, 7102800.0, 7106400.0, 7110000.0, 7113600.0, 7117200.0, 7120800.0, 7124400.0, 7128000.0, 7131600.0, 7135200.0, 7138800.0, 7142400.0, 7146000.0, 7149600.0, 7153200.0, 7156800.0, 7160400.0, 7164000.0, 7167600.0, 7171200.0, 7174800.0, 7178400.0, 7182000.0, 7185600.0, 7189200.0, 7192800.0, 7196400.0, 7200000.0, 7203600.0, 7207200.0, 7210800.0, 7214400.0, 7218000.0, 7221600.0, 7225200.0, 7228800.0, 7232400.0, 7236000.0, 7239600.0, 7243200.0, 7246800.0, 7250400.0, 7254000.0, 7257600.0, 7261200.0, 7264800.0, 7268400.0, 7272000.0, 7275600.0, 7279200.0, 7282800.0, 7286400.0, 7290000.0, 7293600.0, 7297200.0, 7300800.0, 7304400.0, 7308000.0, 7311600.0, 7315200.0, 7318800.0, 7322400.0, 7326000.0, 7329600.0, 7333200.0, 7336800.0, 7340400.0, 7344000.0, 7347600.0, 7351200.0, 7354800.0, 7358400.0, 7362000.0, 7365600.0, 7369200.0, 7372800.0, 7376400.0, 7380000.0, 7383600.0, 7387200.0, 7390800.0, 7394400.0, 7398000.0, 7401600.0, 7405200.0, 7408800.0, 7412400.0, 7416000.0, 7419600.0, 7423200.0, 7426800.0, 7430400.0, 7434000.0, 7437600.0, 7441200.0, 7444800.0, 7448400.0, 7452000.0, 7455600.0, 7459200.0, 7462800.0, 7466400.0, 7470000.0, 7473600.0, 7477200.0, 7480800.0, 7484400.0, 7488000.0, 7491600.0, 7495200.0, 7498800.0, 7502400.0, 7506000.0, 7509600.0, 7513200.0, 7516800.0, 7520400.0, 7524000.0, 7527600.0, 7531200.0, 7534800.0, 7538400.0, 7542000.0, 7545600.0, 7549200.0, 7552800.0, 7556400.0, 7560000.0, 7563600.0, 7567200.0, 7570800.0, 7574400.0, 7578000.0, 7581600.0, 7585200.0, 7588800.0, 7592400.0, 7596000.0, 7599600.0, 7603200.0, 7606800.0, 7610400.0, 7614000.0, 7617600.0, 7621200.0, 7624800.0, 7628400.0, 7632000.0, 7635600.0, 7639200.0, 7642800.0, 7646400.0, 7650000.0, 7653600.0, 7657200.0, 7660800.0, 7664400.0, 7668000.0, 7671600.0, 7675200.0, 7678800.0, 7682400.0, 7686000.0, 7689600.0, 7693200.0, 7696800.0, 7700400.0, 7704000.0, 7707600.0, 7711200.0, 7714800.0, 7718400.0, 7722000.0, 7725600.0, 7729200.0, 7732800.0, 7736400.0, 7740000.0, 7743600.0, 7747200.0, 7750800.0, 7754400.0, 7758000.0, 7761600.0, 7765200.0, 7768800.0, 7772400.0, 7776000.0, 7779600.0, 7783200.0, 7786800.0, 7790400.0, 7794000.0, 7797600.0, 7801200.0, 7804800.0, 7808400.0, 7812000.0, 7815600.0, 7819200.0, 7822800.0, 7826400.0, 7830000.0, 7833600.0, 7837200.0, 7840800.0, 7844400.0, 7848000.0, 7851600.0, 7855200.0, 7858800.0, 7862400.0, 7866000.0, 7869600.0, 7873200.0, 7876800.0, 7880400.0, 7884000.0, 7887600.0, 7891200.0, 7894800.0, 7898400.0, 7902000.0, 7905600.0, 7909200.0, 7912800.0, 7916400.0, 7920000.0, 7923600.0, 7927200.0, 7930800.0, 7934400.0, 7938000.0, 7941600.0, 7945200.0, 7948800.0, 7952400.0, 7956000.0, 7959600.0, 7963200.0, 7966800.0, 7970400.0, 7974000.0, 7977600.0, 7981200.0, 7984800.0, 7988400.0, 7992000.0, 7995600.0, 7999200.0, 8002800.0, 8006400.0, 8010000.0, 8013600.0, 8017200.0, 8020800.0, 8024400.0, 8028000.0, 8031600.0, 8035200.0, 8038800.0, 8042400.0, 8046000.0, 8049600.0, 8053200.0, 8056800.0, 8060400.0, 8064000.0, 8067600.0, 8071200.0, 8074800.0, 8078400.0, 8082000.0, 8085600.0, 8089200.0, 8092800.0, 8096400.0, 8100000.0, 8103600.0, 8107200.0, 8110800.0, 8114400.0, 8118000.0, 8121600.0, 8125200.0, 8128800.0, 8132400.0, 8136000.0, 8139600.0, 8143200.0, 8146800.0, 8150400.0, 8154000.0, 8157600.0, 8161200.0, 8164800.0, 8168400.0, 8172000.0, 8175600.0, 8179200.0, 8182800.0, 8186400.0, 8190000.0, 8193600.0, 8197200.0, 8200800.0, 8204400.0, 8208000.0, 8211600.0, 8215200.0, 8218800.0, 8222400.0, 8226000.0, 8229600.0, 8233200.0, 8236800.0, 8240400.0, 8244000.0, 8247600.0, 8251200.0, 8254800.0, 8258400.0, 8262000.0, 8265600.0, 8269200.0, 8272800.0, 8276400.0, 8280000.0, 8283600.0, 8287200.0, 8290800.0, 8294400.0, 8298000.0, 8301600.0, 8305200.0, 8308800.0, 8312400.0, 8316000.0, 8319600.0, 8323200.0, 8326800.0, 8330400.0, 8334000.0, 8337600.0, 8341200.0, 8344800.0, 8348400.0, 8352000.0, 8355600.0, 8359200.0, 8362800.0, 8366400.0, 8370000.0, 8373600.0, 8377200.0, 8380800.0, 8384400.0, 8388000.0, 8391600.0, 8395200.0, 8398800.0, 8402400.0, 8406000.0, 8409600.0, 8413200.0, 8416800.0, 8420400.0, 8424000.0, 8427600.0, 8431200.0, 8434800.0, 8438400.0, 8442000.0, 8445600.0, 8449200.0, 8452800.0, 8456400.0, 8460000.0, 8463600.0, 8467200.0, 8470800.0, 8474400.0, 8478000.0, 8481600.0, 8485200.0, 8488800.0, 8492400.0, 8496000.0, 8499600.0, 8503200.0, 8506800.0, 8510400.0, 8514000.0, 8517600.0, 8521200.0, 8524800.0, 8528400.0, 8532000.0, 8535600.0, 8539200.0, 8542800.0, 8546400.0, 8550000.0, 8553600.0, 8557200.0, 8560800.0, 8564400.0, 8568000.0, 8571600.0, 8575200.0, 8578800.0, 8582400.0, 8586000.0, 8589600.0, 8593200.0, 8596800.0, 8600400.0, 8604000.0, 8607600.0, 8611200.0, 8614800.0, 8618400.0, 8622000.0, 8625600.0, 8629200.0, 8632800.0, 8636400.0, 8640000.0, 8643600.0, 8647200.0, 8650800.0, 8654400.0, 8658000.0, 8661600.0, 8665200.0, 8668800.0, 8672400.0, 8676000.0, 8679600.0, 8683200.0, 8686800.0, 8690400.0, 8694000.0, 8697600.0, 8701200.0, 8704800.0, 8708400.0, 8712000.0, 8715600.0, 8719200.0, 8722800.0, 8726400.0, 8730000.0, 8733600.0, 8737200.0, 8740800.0, 8744400.0, 8748000.0, 8751600.0, 8755200.0, 8758800.0, 8762400.0, 8766000.0, 8769600.0, 8773200.0, 8776800.0, 8780400.0, 8784000.0, 8787600.0, 8791200.0, 8794800.0, 8798400.0, 8802000.0, 8805600.0, 8809200.0, 8812800.0, 8816400.0, 8820000.0, 8823600.0, 8827200.0, 8830800.0, 8834400.0, 8838000.0, 8841600.0, 8845200.0, 8848800.0, 8852400.0, 8856000.0, 8859600.0, 8863200.0, 8866800.0, 8870400.0, 8874000.0, 8877600.0, 8881200.0, 8884800.0, 8888400.0, 8892000.0, 8895600.0, 8899200.0, 8902800.0, 8906400.0, 8910000.0, 8913600.0, 8917200.0, 8920800.0, 8924400.0, 8928000.0, 8931600.0, 8935200.0, 8938800.0, 8942400.0, 8946000.0, 8949600.0, 8953200.0, 8956800.0, 8960400.0, 8964000.0, 8967600.0, 8971200.0, 8974800.0, 8978400.0, 8982000.0, 8985600.0, 8989200.0, 8992800.0, 8996400.0, 9000000.0, 9003600.0, 9007200.0, 9010800.0, 9014400.0, 9018000.0, 9021600.0, 9025200.0, 9028800.0, 9032400.0, 9036000.0, 9039600.0, 9043200.0, 9046800.0, 9050400.0, 9054000.0, 9057600.0, 9061200.0, 9064800.0, 9068400.0, 9072000.0, 9075600.0, 9079200.0, 9082800.0, 9086400.0, 9090000.0, 9093600.0, 9097200.0, 9100800.0, 9104400.0, 9108000.0, 9111600.0, 9115200.0, 9118800.0, 9122400.0, 9126000.0, 9129600.0, 9133200.0, 9136800.0, 9140400.0, 9144000.0, 9147600.0, 9151200.0, 9154800.0, 9158400.0, 9162000.0, 9165600.0, 9169200.0, 9172800.0, 9176400.0, 9180000.0, 9183600.0, 9187200.0, 9190800.0, 9194400.0, 9198000.0, 9201600.0, 9205200.0, 9208800.0, 9212400.0, 9216000.0, 9219600.0, 9223200.0, 9226800.0, 9230400.0, 9234000.0, 9237600.0, 9241200.0, 9244800.0, 9248400.0, 9252000.0, 9255600.0, 9259200.0, 9262800.0, 9266400.0, 9270000.0, 9273600.0, 9277200.0, 9280800.0, 9284400.0, 9288000.0, 9291600.0, 9295200.0, 9298800.0, 9302400.0, 9306000.0, 9309600.0, 9313200.0, 9316800.0, 9320400.0, 9324000.0, 9327600.0, 9331200.0, 9334800.0, 9338400.0, 9342000.0, 9345600.0, 9349200.0, 9352800.0, 9356400.0, 9360000.0, 9363600.0, 9367200.0, 9370800.0, 9374400.0, 9378000.0, 9381600.0, 9385200.0, 9388800.0, 9392400.0, 9396000.0, 9399600.0, 9403200.0, 9406800.0, 9410400.0, 9414000.0, 9417600.0, 9421200.0, 9424800.0, 9428400.0, 9432000.0, 9435600.0, 9439200.0, 9442800.0, 9446400.0, 9450000.0, 9453600.0, 9457200.0, 9460800.0, 9464400.0, 9468000.0, 9471600.0, 9475200.0, 9478800.0, 9482400.0, 9486000.0, 9489600.0, 9493200.0, 9496800.0, 9500400.0, 9504000.0, 9507600.0, 9511200.0, 9514800.0, 9518400.0, 9522000.0, 9525600.0, 9529200.0, 9532800.0, 9536400.0, 9540000.0, 9543600.0, 9547200.0, 9550800.0, 9554400.0, 9558000.0, 9561600.0, 9565200.0, 9568800.0, 9572400.0, 9576000.0, 9579600.0, 9583200.0, 9586800.0, 9590400.0, 9594000.0, 9597600.0, 9601200.0, 9604800.0, 9608400.0, 9612000.0, 9615600.0, 9619200.0, 9622800.0, 9626400.0, 9630000.0, 9633600.0, 9637200.0, 9640800.0, 9644400.0, 9648000.0, 9651600.0, 9655200.0, 9658800.0, 9662400.0, 9666000.0, 9669600.0, 9673200.0, 9676800.0, 9680400.0, 9684000.0, 9687600.0, 9691200.0, 9694800.0, 9698400.0, 9702000.0, 9705600.0, 9709200.0, 9712800.0, 9716400.0, 9720000.0, 9723600.0, 9727200.0, 9730800.0, 9734400.0, 9738000.0, 9741600.0, 9745200.0, 9748800.0, 9752400.0, 9756000.0, 9759600.0, 9763200.0, 9766800.0, 9770400.0, 9774000.0, 9777600.0, 9781200.0, 9784800.0, 9788400.0, 9792000.0, 9795600.0, 9799200.0, 9802800.0, 9806400.0, 9810000.0, 9813600.0, 9817200.0, 9820800.0, 9824400.0, 9828000.0, 9831600.0, 9835200.0, 9838800.0, 9842400.0, 9846000.0, 9849600.0, 9853200.0, 9856800.0, 9860400.0, 9864000.0, 9867600.0, 9871200.0, 9874800.0, 9878400.0, 9882000.0, 9885600.0, 9889200.0, 9892800.0, 9896400.0, 9900000.0, 9903600.0, 9907200.0, 9910800.0, 9914400.0, 9918000.0, 9921600.0, 9925200.0, 9928800.0, 9932400.0, 9936000.0, 9939600.0, 9943200.0, 9946800.0, 9950400.0, 9954000.0, 9957600.0, 9961200.0, 9964800.0, 9968400.0, 9972000.0, 9975600.0, 9979200.0, 9982800.0, 9986400.0, 9990000.0, 9993600.0, 9997200.0, 10000800.0, 10004400.0, 10008000.0, 10011600.0, 10015200.0, 10018800.0, 10022400.0, 10026000.0, 10029600.0, 10033200.0, 10036800.0, 10040400.0, 10044000.0, 10047600.0, 10051200.0, 10054800.0, 10058400.0, 10062000.0, 10065600.0, 10069200.0, 10072800.0, 10076400.0, 10080000.0, 10083600.0, 10087200.0, 10090800.0, 10094400.0, 10098000.0, 10101600.0, 10105200.0, 10108800.0, 10112400.0, 10116000.0, 10119600.0, 10123200.0, 10126800.0, 10130400.0, 10134000.0, 10137600.0, 10141200.0, 10144800.0, 10148400.0, 10152000.0, 10155600.0, 10159200.0, 10162800.0, 10166400.0, 10170000.0, 10173600.0, 10177200.0, 10180800.0, 10184400.0, 10188000.0, 10191600.0, 10195200.0, 10198800.0, 10202400.0, 10206000.0, 10209600.0, 10213200.0, 10216800.0, 10220400.0, 10224000.0, 10227600.0, 10231200.0, 10234800.0, 10238400.0, 10242000.0, 10245600.0, 10249200.0, 10252800.0, 10256400.0, 10260000.0, 10263600.0, 10267200.0, 10270800.0, 10274400.0, 10278000.0, 10281600.0, 10285200.0, 10288800.0, 10292400.0, 10296000.0, 10299600.0, 10303200.0, 10306800.0, 10310400.0, 10314000.0, 10317600.0, 10321200.0, 10324800.0, 10328400.0, 10332000.0, 10335600.0, 10339200.0, 10342800.0, 10346400.0, 10350000.0, 10353600.0, 10357200.0, 10360800.0, 10364400.0, 10368000.0, 10371600.0, 10375200.0, 10378800.0, 10382400.0, 10386000.0, 10389600.0, 10393200.0, 10396800.0, 10400400.0, 10404000.0, 10407600.0, 10411200.0, 10414800.0, 10418400.0, 10422000.0, 10425600.0, 10429200.0, 10432800.0, 10436400.0, 10440000.0, 10443600.0, 10447200.0, 10450800.0, 10454400.0, 10458000.0, 10461600.0, 10465200.0, 10468800.0, 10472400.0, 10476000.0, 10479600.0, 10483200.0, 10486800.0, 10490400.0, 10494000.0, 10497600.0, 10501200.0, 10504800.0, 10508400.0, 10512000.0, 10515600.0, 10519200.0, 10522800.0, 10526400.0, 10530000.0, 10533600.0, 10537200.0, 10540800.0, 10544400.0, 10548000.0, 10551600.0, 10555200.0, 10558800.0, 10562400.0, 10566000.0, 10569600.0, 10573200.0, 10576800.0, 10580400.0, 10584000.0, 10587600.0, 10591200.0, 10594800.0, 10598400.0, 10602000.0, 10605600.0, 10609200.0, 10612800.0, 10616400.0, 10620000.0, 10623600.0, 10627200.0, 10630800.0, 10634400.0, 10638000.0, 10641600.0, 10645200.0, 10648800.0, 10652400.0, 10656000.0, 10659600.0, 10663200.0, 10666800.0, 10670400.0, 10674000.0, 10677600.0, 10681200.0, 10684800.0, 10688400.0, 10692000.0, 10695600.0, 10699200.0, 10702800.0, 10706400.0, 10710000.0, 10713600.0, 10717200.0, 10720800.0, 10724400.0, 10728000.0, 10731600.0, 10735200.0, 10738800.0, 10742400.0, 10746000.0, 10749600.0, 10753200.0, 10756800.0, 10760400.0, 10764000.0, 10767600.0, 10771200.0, 10774800.0, 10778400.0, 10782000.0, 10785600.0, 10789200.0, 10792800.0, 10796400.0, 10800000.0, 10803600.0, 10807200.0, 10810800.0, 10814400.0, 10818000.0, 10821600.0, 10825200.0, 10828800.0, 10832400.0, 10836000.0, 10839600.0, 10843200.0, 10846800.0, 10850400.0, 10854000.0, 10857600.0, 10861200.0, 10864800.0, 10868400.0, 10872000.0, 10875600.0, 10879200.0, 10882800.0, 10886400.0, 10890000.0, 10893600.0, 10897200.0, 10900800.0, 10904400.0, 10908000.0, 10911600.0, 10915200.0, 10918800.0, 10922400.0, 10926000.0, 10929600.0, 10933200.0, 10936800.0, 10940400.0, 10944000.0, 10947600.0, 10951200.0, 10954800.0, 10958400.0, 10962000.0, 10965600.0, 10969200.0, 10972800.0, 10976400.0, 10980000.0, 10983600.0, 10987200.0, 10990800.0, 10994400.0, 10998000.0, 11001600.0, 11005200.0, 11008800.0, 11012400.0, 11016000.0, 11019600.0, 11023200.0, 11026800.0, 11030400.0, 11034000.0, 11037600.0, 11041200.0, 11044800.0, 11048400.0, 11052000.0, 11055600.0, 11059200.0, 11062800.0, 11066400.0, 11070000.0, 11073600.0, 11077200.0, 11080800.0, 11084400.0, 11088000.0, 11091600.0, 11095200.0, 11098800.0, 11102400.0, 11106000.0, 11109600.0, 11113200.0, 11116800.0, 11120400.0, 11124000.0, 11127600.0, 11131200.0, 11134800.0, 11138400.0, 11142000.0, 11145600.0, 11149200.0, 11152800.0, 11156400.0, 11160000.0, 11163600.0, 11167200.0, 11170800.0, 11174400.0, 11178000.0, 11181600.0, 11185200.0, 11188800.0, 11192400.0, 11196000.0, 11199600.0, 11203200.0, 11206800.0, 11210400.0, 11214000.0, 11217600.0, 11221200.0, 11224800.0, 11228400.0, 11232000.0, 11235600.0, 11239200.0, 11242800.0, 11246400.0, 11250000.0, 11253600.0, 11257200.0, 11260800.0, 11264400.0, 11268000.0, 11271600.0, 11275200.0, 11278800.0, 11282400.0, 11286000.0, 11289600.0, 11293200.0, 11296800.0, 11300400.0, 11304000.0, 11307600.0, 11311200.0, 11314800.0, 11318400.0, 11322000.0, 11325600.0, 11329200.0, 11332800.0, 11336400.0, 11340000.0, 11343600.0, 11347200.0, 11350800.0, 11354400.0, 11358000.0, 11361600.0, 11365200.0, 11368800.0, 11372400.0, 11376000.0, 11379600.0, 11383200.0, 11386800.0, 11390400.0, 11394000.0, 11397600.0, 11401200.0, 11404800.0, 11408400.0, 11412000.0, 11415600.0, 11419200.0, 11422800.0, 11426400.0, 11430000.0, 11433600.0, 11437200.0, 11440800.0, 11444400.0, 11448000.0, 11451600.0, 11455200.0, 11458800.0, 11462400.0, 11466000.0, 11469600.0, 11473200.0, 11476800.0, 11480400.0, 11484000.0, 11487600.0, 11491200.0, 11494800.0, 11498400.0, 11502000.0, 11505600.0, 11509200.0, 11512800.0, 11516400.0, 11520000.0, 11523600.0, 11527200.0, 11530800.0, 11534400.0, 11538000.0, 11541600.0, 11545200.0, 11548800.0, 11552400.0, 11556000.0, 11559600.0, 11563200.0, 11566800.0, 11570400.0, 11574000.0, 11577600.0, 11581200.0, 11584800.0, 11588400.0, 11592000.0, 11595600.0, 11599200.0, 11602800.0, 11606400.0, 11610000.0, 11613600.0, 11617200.0, 11620800.0, 11624400.0, 11628000.0, 11631600.0, 11635200.0, 11638800.0, 11642400.0, 11646000.0, 11649600.0, 11653200.0, 11656800.0, 11660400.0, 11664000.0, 11667600.0, 11671200.0, 11674800.0, 11678400.0, 11682000.0, 11685600.0, 11689200.0, 11692800.0, 11696400.0, 11700000.0, 11703600.0, 11707200.0, 11710800.0, 11714400.0, 11718000.0, 11721600.0, 11725200.0, 11728800.0, 11732400.0, 11736000.0, 11739600.0, 11743200.0, 11746800.0, 11750400.0, 11754000.0, 11757600.0, 11761200.0, 11764800.0, 11768400.0, 11772000.0, 11775600.0, 11779200.0, 11782800.0, 11786400.0, 11790000.0, 11793600.0, 11797200.0, 11800800.0, 11804400.0, 11808000.0, 11811600.0, 11815200.0, 11818800.0, 11822400.0, 11826000.0, 11829600.0, 11833200.0, 11836800.0, 11840400.0, 11844000.0, 11847600.0, 11851200.0, 11854800.0, 11858400.0, 11862000.0, 11865600.0, 11869200.0, 11872800.0, 11876400.0, 11880000.0, 11883600.0, 11887200.0, 11890800.0, 11894400.0, 11898000.0, 11901600.0, 11905200.0, 11908800.0, 11912400.0, 11916000.0, 11919600.0, 11923200.0, 11926800.0, 11930400.0, 11934000.0, 11937600.0, 11941200.0, 11944800.0, 11948400.0, 11952000.0, 11955600.0, 11959200.0, 11962800.0, 11966400.0, 11970000.0, 11973600.0, 11977200.0, 11980800.0, 11984400.0, 11988000.0, 11991600.0, 11995200.0, 11998800.0, 12002400.0, 12006000.0, 12009600.0, 12013200.0, 12016800.0, 12020400.0, 12024000.0, 12027600.0, 12031200.0, 12034800.0, 12038400.0, 12042000.0, 12045600.0, 12049200.0, 12052800.0, 12056400.0, 12060000.0, 12063600.0, 12067200.0, 12070800.0, 12074400.0, 12078000.0, 12081600.0, 12085200.0, 12088800.0, 12092400.0, 12096000.0, 12099600.0, 12103200.0, 12106800.0, 12110400.0, 12114000.0, 12117600.0, 12121200.0, 12124800.0, 12128400.0, 12132000.0, 12135600.0, 12139200.0, 12142800.0, 12146400.0, 12150000.0, 12153600.0, 12157200.0, 12160800.0, 12164400.0, 12168000.0, 12171600.0, 12175200.0, 12178800.0, 12182400.0, 12186000.0, 12189600.0, 12193200.0, 12196800.0, 12200400.0, 12204000.0, 12207600.0, 12211200.0, 12214800.0, 12218400.0, 12222000.0, 12225600.0, 12229200.0, 12232800.0, 12236400.0, 12240000.0, 12243600.0, 12247200.0, 12250800.0, 12254400.0, 12258000.0, 12261600.0, 12265200.0, 12268800.0, 12272400.0, 12276000.0, 12279600.0, 12283200.0, 12286800.0, 12290400.0, 12294000.0, 12297600.0, 12301200.0, 12304800.0, 12308400.0, 12312000.0, 12315600.0, 12319200.0, 12322800.0, 12326400.0, 12330000.0, 12333600.0, 12337200.0, 12340800.0, 12344400.0, 12348000.0, 12351600.0, 12355200.0, 12358800.0, 12362400.0, 12366000.0, 12369600.0, 12373200.0, 12376800.0, 12380400.0, 12384000.0, 12387600.0, 12391200.0, 12394800.0, 12398400.0, 12402000.0, 12405600.0, 12409200.0, 12412800.0, 12416400.0, 12420000.0, 12423600.0, 12427200.0, 12430800.0, 12434400.0, 12438000.0, 12441600.0, 12445200.0, 12448800.0, 12452400.0, 12456000.0, 12459600.0, 12463200.0, 12466800.0, 12470400.0, 12474000.0, 12477600.0, 12481200.0, 12484800.0, 12488400.0, 12492000.0, 12495600.0, 12499200.0, 12502800.0, 12506400.0, 12510000.0, 12513600.0, 12517200.0, 12520800.0, 12524400.0, 12528000.0, 12531600.0, 12535200.0, 12538800.0, 12542400.0, 12546000.0, 12549600.0, 12553200.0, 12556800.0, 12560400.0, 12564000.0, 12567600.0, 12571200.0, 12574800.0, 12578400.0, 12582000.0, 12585600.0, 12589200.0, 12592800.0, 12596400.0, 12600000.0, 12603600.0, 12607200.0, 12610800.0, 12614400.0, 12618000.0, 12621600.0, 12625200.0, 12628800.0, 12632400.0, 12636000.0, 12639600.0, 12643200.0, 12646800.0, 12650400.0, 12654000.0, 12657600.0, 12661200.0, 12664800.0, 12668400.0, 12672000.0, 12675600.0, 12679200.0, 12682800.0, 12686400.0, 12690000.0, 12693600.0, 12697200.0, 12700800.0, 12704400.0, 12708000.0, 12711600.0, 12715200.0, 12718800.0, 12722400.0, 12726000.0, 12729600.0, 12733200.0, 12736800.0, 12740400.0, 12744000.0, 12747600.0, 12751200.0, 12754800.0, 12758400.0, 12762000.0, 12765600.0, 12769200.0, 12772800.0, 12776400.0, 12780000.0, 12783600.0, 12787200.0, 12790800.0, 12794400.0, 12798000.0, 12801600.0, 12805200.0, 12808800.0, 12812400.0, 12816000.0, 12819600.0, 12823200.0, 12826800.0, 12830400.0, 12834000.0, 12837600.0, 12841200.0, 12844800.0, 12848400.0, 12852000.0, 12855600.0, 12859200.0, 12862800.0, 12866400.0, 12870000.0, 12873600.0, 12877200.0, 12880800.0, 12884400.0, 12888000.0, 12891600.0, 12895200.0, 12898800.0, 12902400.0, 12906000.0, 12909600.0, 12913200.0, 12916800.0, 12920400.0, 12924000.0, 12927600.0, 12931200.0, 12934800.0, 12938400.0, 12942000.0, 12945600.0, 12949200.0, 12952800.0, 12956400.0, 12960000.0, 12963600.0, 12967200.0, 12970800.0, 12974400.0, 12978000.0, 12981600.0, 12985200.0, 12988800.0, 12992400.0, 12996000.0, 12999600.0, 13003200.0, 13006800.0, 13010400.0, 13014000.0, 13017600.0, 13021200.0, 13024800.0, 13028400.0, 13032000.0, 13035600.0, 13039200.0, 13042800.0, 13046400.0, 13050000.0, 13053600.0, 13057200.0, 13060800.0, 13064400.0, 13068000.0, 13071600.0, 13075200.0, 13078800.0, 13082400.0, 13086000.0, 13089600.0, 13093200.0, 13096800.0, 13100400.0, 13104000.0, 13107600.0, 13111200.0, 13114800.0, 13118400.0, 13122000.0, 13125600.0, 13129200.0, 13132800.0, 13136400.0, 13140000.0, 13143600.0, 13147200.0, 13150800.0, 13154400.0, 13158000.0, 13161600.0, 13165200.0, 13168800.0, 13172400.0, 13176000.0, 13179600.0, 13183200.0, 13186800.0, 13190400.0, 13194000.0, 13197600.0, 13201200.0, 13204800.0, 13208400.0, 13212000.0, 13215600.0, 13219200.0, 13222800.0, 13226400.0, 13230000.0, 13233600.0, 13237200.0, 13240800.0, 13244400.0, 13248000.0, 13251600.0, 13255200.0, 13258800.0, 13262400.0, 13266000.0, 13269600.0, 13273200.0, 13276800.0, 13280400.0, 13284000.0, 13287600.0, 13291200.0, 13294800.0, 13298400.0, 13302000.0, 13305600.0, 13309200.0, 13312800.0, 13316400.0, 13320000.0, 13323600.0, 13327200.0, 13330800.0, 13334400.0, 13338000.0, 13341600.0, 13345200.0, 13348800.0, 13352400.0, 13356000.0, 13359600.0, 13363200.0, 13366800.0, 13370400.0, 13374000.0, 13377600.0, 13381200.0, 13384800.0, 13388400.0, 13392000.0, 13395600.0, 13399200.0, 13402800.0, 13406400.0, 13410000.0, 13413600.0, 13417200.0, 13420800.0, 13424400.0, 13428000.0, 13431600.0, 13435200.0, 13438800.0, 13442400.0, 13446000.0, 13449600.0, 13453200.0, 13456800.0, 13460400.0, 13464000.0, 13467600.0, 13471200.0, 13474800.0, 13478400.0, 13482000.0, 13485600.0, 13489200.0, 13492800.0, 13496400.0, 13500000.0, 13503600.0, 13507200.0, 13510800.0, 13514400.0, 13518000.0, 13521600.0, 13525200.0, 13528800.0, 13532400.0, 13536000.0, 13539600.0, 13543200.0, 13546800.0, 13550400.0, 13554000.0, 13557600.0, 13561200.0, 13564800.0, 13568400.0, 13572000.0, 13575600.0, 13579200.0, 13582800.0, 13586400.0, 13590000.0, 13593600.0, 13597200.0, 13600800.0, 13604400.0, 13608000.0, 13611600.0, 13615200.0, 13618800.0, 13622400.0, 13626000.0, 13629600.0, 13633200.0, 13636800.0, 13640400.0, 13644000.0, 13647600.0, 13651200.0, 13654800.0, 13658400.0, 13662000.0, 13665600.0, 13669200.0, 13672800.0, 13676400.0, 13680000.0, 13683600.0, 13687200.0, 13690800.0, 13694400.0, 13698000.0, 13701600.0, 13705200.0, 13708800.0, 13712400.0, 13716000.0, 13719600.0, 13723200.0, 13726800.0, 13730400.0, 13734000.0, 13737600.0, 13741200.0, 13744800.0, 13748400.0, 13752000.0, 13755600.0, 13759200.0, 13762800.0, 13766400.0, 13770000.0, 13773600.0, 13777200.0, 13780800.0, 13784400.0, 13788000.0, 13791600.0, 13795200.0, 13798800.0, 13802400.0, 13806000.0, 13809600.0, 13813200.0, 13816800.0, 13820400.0, 13824000.0, 13827600.0, 13831200.0, 13834800.0, 13838400.0, 13842000.0, 13845600.0, 13849200.0, 13852800.0, 13856400.0, 13860000.0, 13863600.0, 13867200.0, 13870800.0, 13874400.0, 13878000.0, 13881600.0, 13885200.0, 13888800.0, 13892400.0, 13896000.0, 13899600.0, 13903200.0, 13906800.0, 13910400.0, 13914000.0, 13917600.0, 13921200.0, 13924800.0, 13928400.0, 13932000.0, 13935600.0, 13939200.0, 13942800.0, 13946400.0, 13950000.0, 13953600.0, 13957200.0, 13960800.0, 13964400.0, 13968000.0, 13971600.0, 13975200.0, 13978800.0, 13982400.0, 13986000.0, 13989600.0, 13993200.0, 13996800.0, 14000400.0, 14004000.0, 14007600.0, 14011200.0, 14014800.0, 14018400.0, 14022000.0, 14025600.0, 14029200.0, 14032800.0, 14036400.0, 14040000.0, 14043600.0, 14047200.0, 14050800.0, 14054400.0, 14058000.0, 14061600.0, 14065200.0, 14068800.0, 14072400.0, 14076000.0, 14079600.0, 14083200.0, 14086800.0, 14090400.0, 14094000.0, 14097600.0, 14101200.0, 14104800.0, 14108400.0, 14112000.0, 14115600.0, 14119200.0, 14122800.0, 14126400.0, 14130000.0, 14133600.0, 14137200.0, 14140800.0, 14144400.0, 14148000.0, 14151600.0, 14155200.0, 14158800.0, 14162400.0, 14166000.0, 14169600.0, 14173200.0, 14176800.0, 14180400.0, 14184000.0, 14187600.0, 14191200.0, 14194800.0, 14198400.0, 14202000.0, 14205600.0, 14209200.0, 14212800.0, 14216400.0, 14220000.0, 14223600.0, 14227200.0, 14230800.0, 14234400.0, 14238000.0, 14241600.0, 14245200.0, 14248800.0, 14252400.0, 14256000.0, 14259600.0, 14263200.0, 14266800.0, 14270400.0, 14274000.0, 14277600.0, 14281200.0, 14284800.0, 14288400.0, 14292000.0, 14295600.0, 14299200.0, 14302800.0, 14306400.0, 14310000.0, 14313600.0, 14317200.0, 14320800.0, 14324400.0, 14328000.0, 14331600.0, 14335200.0, 14338800.0, 14342400.0, 14346000.0, 14349600.0, 14353200.0, 14356800.0, 14360400.0, 14364000.0, 14367600.0, 14371200.0, 14374800.0, 14378400.0, 14382000.0, 14385600.0, 14389200.0, 14392800.0, 14396400.0, 14400000.0, 14403600.0, 14407200.0, 14410800.0, 14414400.0, 14418000.0, 14421600.0, 14425200.0, 14428800.0, 14432400.0, 14436000.0, 14439600.0, 14443200.0, 14446800.0, 14450400.0, 14454000.0, 14457600.0, 14461200.0, 14464800.0, 14468400.0, 14472000.0, 14475600.0, 14479200.0, 14482800.0, 14486400.0, 14490000.0, 14493600.0, 14497200.0, 14500800.0, 14504400.0, 14508000.0, 14511600.0, 14515200.0, 14518800.0, 14522400.0, 14526000.0, 14529600.0, 14533200.0, 14536800.0, 14540400.0, 14544000.0, 14547600.0, 14551200.0, 14554800.0, 14558400.0, 14562000.0, 14565600.0, 14569200.0, 14572800.0, 14576400.0, 14580000.0, 14583600.0, 14587200.0, 14590800.0, 14594400.0, 14598000.0, 14601600.0, 14605200.0, 14608800.0, 14612400.0, 14616000.0, 14619600.0, 14623200.0, 14626800.0, 14630400.0, 14634000.0, 14637600.0, 14641200.0, 14644800.0, 14648400.0, 14652000.0, 14655600.0, 14659200.0, 14662800.0, 14666400.0, 14670000.0, 14673600.0, 14677200.0, 14680800.0, 14684400.0, 14688000.0, 14691600.0, 14695200.0, 14698800.0, 14702400.0, 14706000.0, 14709600.0, 14713200.0, 14716800.0, 14720400.0, 14724000.0, 14727600.0, 14731200.0, 14734800.0, 14738400.0, 14742000.0, 14745600.0, 14749200.0, 14752800.0, 14756400.0, 14760000.0, 14763600.0, 14767200.0, 14770800.0, 14774400.0, 14778000.0, 14781600.0, 14785200.0, 14788800.0, 14792400.0, 14796000.0, 14799600.0, 14803200.0, 14806800.0, 14810400.0, 14814000.0, 14817600.0, 14821200.0, 14824800.0, 14828400.0, 14832000.0, 14835600.0, 14839200.0, 14842800.0, 14846400.0, 14850000.0, 14853600.0, 14857200.0, 14860800.0, 14864400.0, 14868000.0, 14871600.0, 14875200.0, 14878800.0, 14882400.0, 14886000.0, 14889600.0, 14893200.0, 14896800.0, 14900400.0, 14904000.0, 14907600.0, 14911200.0, 14914800.0, 14918400.0, 14922000.0, 14925600.0, 14929200.0, 14932800.0, 14936400.0, 14940000.0, 14943600.0, 14947200.0, 14950800.0, 14954400.0, 14958000.0, 14961600.0, 14965200.0, 14968800.0, 14972400.0, 14976000.0, 14979600.0, 14983200.0, 14986800.0, 14990400.0, 14994000.0, 14997600.0, 15001200.0, 15004800.0, 15008400.0, 15012000.0, 15015600.0, 15019200.0, 15022800.0, 15026400.0, 15030000.0, 15033600.0, 15037200.0, 15040800.0, 15044400.0, 15048000.0, 15051600.0, 15055200.0, 15058800.0, 15062400.0, 15066000.0, 15069600.0, 15073200.0, 15076800.0, 15080400.0, 15084000.0, 15087600.0, 15091200.0, 15094800.0, 15098400.0, 15102000.0, 15105600.0, 15109200.0, 15112800.0, 15116400.0, 15120000.0, 15123600.0, 15127200.0, 15130800.0, 15134400.0, 15138000.0, 15141600.0, 15145200.0, 15148800.0, 15152400.0, 15156000.0, 15159600.0, 15163200.0, 15166800.0, 15170400.0, 15174000.0, 15177600.0, 15181200.0, 15184800.0, 15188400.0, 15192000.0, 15195600.0, 15199200.0, 15202800.0, 15206400.0, 15210000.0, 15213600.0, 15217200.0, 15220800.0, 15224400.0, 15228000.0, 15231600.0, 15235200.0, 15238800.0, 15242400.0, 15246000.0, 15249600.0, 15253200.0, 15256800.0, 15260400.0, 15264000.0, 15267600.0, 15271200.0, 15274800.0, 15278400.0, 15282000.0, 15285600.0, 15289200.0, 15292800.0, 15296400.0, 15300000.0, 15303600.0, 15307200.0, 15310800.0, 15314400.0, 15318000.0, 15321600.0, 15325200.0, 15328800.0, 15332400.0, 15336000.0, 15339600.0, 15343200.0, 15346800.0, 15350400.0, 15354000.0, 15357600.0, 15361200.0, 15364800.0, 15368400.0, 15372000.0, 15375600.0, 15379200.0, 15382800.0, 15386400.0, 15390000.0, 15393600.0, 15397200.0, 15400800.0, 15404400.0, 15408000.0, 15411600.0, 15415200.0, 15418800.0, 15422400.0, 15426000.0, 15429600.0, 15433200.0, 15436800.0, 15440400.0, 15444000.0, 15447600.0, 15451200.0, 15454800.0, 15458400.0, 15462000.0, 15465600.0, 15469200.0, 15472800.0, 15476400.0, 15480000.0, 15483600.0, 15487200.0, 15490800.0, 15494400.0, 15498000.0, 15501600.0, 15505200.0, 15508800.0, 15512400.0, 15516000.0, 15519600.0, 15523200.0, 15526800.0, 15530400.0, 15534000.0, 15537600.0, 15541200.0, 15544800.0, 15548400.0, 15552000.0, 15555600.0, 15559200.0, 15562800.0, 15566400.0, 15570000.0, 15573600.0, 15577200.0, 15580800.0, 15584400.0, 15588000.0, 15591600.0, 15595200.0, 15598800.0, 15602400.0, 15606000.0, 15609600.0, 15613200.0, 15616800.0, 15620400.0, 15624000.0, 15627600.0, 15631200.0, 15634800.0, 15638400.0, 15642000.0, 15645600.0, 15649200.0, 15652800.0, 15656400.0, 15660000.0, 15663600.0, 15667200.0, 15670800.0, 15674400.0, 15678000.0, 15681600.0, 15685200.0, 15688800.0, 15692400.0, 15696000.0, 15699600.0, 15703200.0, 15706800.0, 15710400.0, 15714000.0, 15717600.0, 15721200.0, 15724800.0, 15728400.0, 15732000.0, 15735600.0, 15739200.0, 15742800.0, 15746400.0, 15750000.0, 15753600.0, 15757200.0, 15760800.0, 15764400.0, 15768000.0, 15771600.0, 15775200.0, 15778800.0, 15782400.0, 15786000.0, 15789600.0, 15793200.0, 15796800.0, 15800400.0, 15804000.0, 15807600.0, 15811200.0, 15814800.0, 15818400.0, 15822000.0, 15825600.0, 15829200.0, 15832800.0, 15836400.0, 15840000.0, 15843600.0, 15847200.0, 15850800.0, 15854400.0, 15858000.0, 15861600.0, 15865200.0, 15868800.0, 15872400.0, 15876000.0, 15879600.0, 15883200.0, 15886800.0, 15890400.0, 15894000.0, 15897600.0, 15901200.0, 15904800.0, 15908400.0, 15912000.0, 15915600.0, 15919200.0, 15922800.0, 15926400.0, 15930000.0, 15933600.0, 15937200.0, 15940800.0, 15944400.0, 15948000.0, 15951600.0, 15955200.0, 15958800.0, 15962400.0, 15966000.0, 15969600.0, 15973200.0, 15976800.0, 15980400.0, 15984000.0, 15987600.0, 15991200.0, 15994800.0, 15998400.0, 16002000.0, 16005600.0, 16009200.0, 16012800.0, 16016400.0, 16020000.0, 16023600.0, 16027200.0, 16030800.0, 16034400.0, 16038000.0, 16041600.0, 16045200.0, 16048800.0, 16052400.0, 16056000.0, 16059600.0, 16063200.0, 16066800.0, 16070400.0, 16074000.0, 16077600.0, 16081200.0, 16084800.0, 16088400.0, 16092000.0, 16095600.0, 16099200.0, 16102800.0, 16106400.0, 16110000.0, 16113600.0, 16117200.0, 16120800.0, 16124400.0, 16128000.0, 16131600.0, 16135200.0, 16138800.0, 16142400.0, 16146000.0, 16149600.0, 16153200.0, 16156800.0, 16160400.0, 16164000.0, 16167600.0, 16171200.0, 16174800.0, 16178400.0, 16182000.0, 16185600.0, 16189200.0, 16192800.0, 16196400.0, 16200000.0, 16203600.0, 16207200.0, 16210800.0, 16214400.0, 16218000.0, 16221600.0, 16225200.0, 16228800.0, 16232400.0, 16236000.0, 16239600.0, 16243200.0, 16246800.0, 16250400.0, 16254000.0, 16257600.0, 16261200.0, 16264800.0, 16268400.0, 16272000.0, 16275600.0, 16279200.0, 16282800.0, 16286400.0, 16290000.0, 16293600.0, 16297200.0, 16300800.0, 16304400.0, 16308000.0, 16311600.0, 16315200.0, 16318800.0, 16322400.0, 16326000.0, 16329600.0, 16333200.0, 16336800.0, 16340400.0, 16344000.0, 16347600.0, 16351200.0, 16354800.0, 16358400.0, 16362000.0, 16365600.0, 16369200.0, 16372800.0, 16376400.0, 16380000.0, 16383600.0, 16387200.0, 16390800.0, 16394400.0, 16398000.0, 16401600.0, 16405200.0, 16408800.0, 16412400.0, 16416000.0, 16419600.0, 16423200.0, 16426800.0, 16430400.0, 16434000.0, 16437600.0, 16441200.0, 16444800.0, 16448400.0, 16452000.0, 16455600.0, 16459200.0, 16462800.0, 16466400.0, 16470000.0, 16473600.0, 16477200.0, 16480800.0, 16484400.0, 16488000.0, 16491600.0, 16495200.0, 16498800.0, 16502400.0, 16506000.0, 16509600.0, 16513200.0, 16516800.0, 16520400.0, 16524000.0, 16527600.0, 16531200.0, 16534800.0, 16538400.0, 16542000.0, 16545600.0, 16549200.0, 16552800.0, 16556400.0, 16560000.0, 16563600.0, 16567200.0, 16570800.0, 16574400.0, 16578000.0, 16581600.0, 16585200.0, 16588800.0, 16592400.0, 16596000.0, 16599600.0, 16603200.0, 16606800.0, 16610400.0, 16614000.0, 16617600.0, 16621200.0, 16624800.0, 16628400.0, 16632000.0, 16635600.0, 16639200.0, 16642800.0, 16646400.0, 16650000.0, 16653600.0, 16657200.0, 16660800.0, 16664400.0, 16668000.0, 16671600.0, 16675200.0, 16678800.0, 16682400.0, 16686000.0, 16689600.0, 16693200.0, 16696800.0, 16700400.0, 16704000.0, 16707600.0, 16711200.0, 16714800.0, 16718400.0, 16722000.0, 16725600.0, 16729200.0, 16732800.0, 16736400.0, 16740000.0, 16743600.0, 16747200.0, 16750800.0, 16754400.0, 16758000.0, 16761600.0, 16765200.0, 16768800.0, 16772400.0, 16776000.0, 16779600.0, 16783200.0, 16786800.0, 16790400.0, 16794000.0, 16797600.0, 16801200.0, 16804800.0, 16808400.0, 16812000.0, 16815600.0, 16819200.0, 16822800.0, 16826400.0, 16830000.0, 16833600.0, 16837200.0, 16840800.0, 16844400.0, 16848000.0, 16851600.0, 16855200.0, 16858800.0, 16862400.0, 16866000.0, 16869600.0, 16873200.0, 16876800.0, 16880400.0, 16884000.0, 16887600.0, 16891200.0, 16894800.0, 16898400.0, 16902000.0, 16905600.0, 16909200.0, 16912800.0, 16916400.0, 16920000.0, 16923600.0, 16927200.0, 16930800.0, 16934400.0, 16938000.0, 16941600.0, 16945200.0, 16948800.0, 16952400.0, 16956000.0, 16959600.0, 16963200.0, 16966800.0, 16970400.0, 16974000.0, 16977600.0, 16981200.0, 16984800.0, 16988400.0, 16992000.0, 16995600.0, 16999200.0, 17002800.0, 17006400.0, 17010000.0, 17013600.0, 17017200.0, 17020800.0, 17024400.0, 17028000.0, 17031600.0, 17035200.0, 17038800.0, 17042400.0, 17046000.0, 17049600.0, 17053200.0, 17056800.0, 17060400.0, 17064000.0, 17067600.0, 17071200.0, 17074800.0, 17078400.0, 17082000.0, 17085600.0, 17089200.0, 17092800.0, 17096400.0, 17100000.0, 17103600.0, 17107200.0, 17110800.0, 17114400.0, 17118000.0, 17121600.0, 17125200.0, 17128800.0, 17132400.0, 17136000.0, 17139600.0, 17143200.0, 17146800.0, 17150400.0, 17154000.0, 17157600.0, 17161200.0, 17164800.0, 17168400.0, 17172000.0, 17175600.0, 17179200.0, 17182800.0, 17186400.0, 17190000.0, 17193600.0, 17197200.0, 17200800.0, 17204400.0, 17208000.0, 17211600.0, 17215200.0, 17218800.0, 17222400.0, 17226000.0, 17229600.0, 17233200.0, 17236800.0, 17240400.0, 17244000.0, 17247600.0, 17251200.0, 17254800.0, 17258400.0, 17262000.0, 17265600.0, 17269200.0, 17272800.0, 17276400.0, 17280000.0, 17283600.0, 17287200.0, 17290800.0, 17294400.0, 17298000.0, 17301600.0, 17305200.0, 17308800.0, 17312400.0, 17316000.0, 17319600.0, 17323200.0, 17326800.0, 17330400.0, 17334000.0, 17337600.0, 17341200.0, 17344800.0, 17348400.0, 17352000.0, 17355600.0, 17359200.0, 17362800.0, 17366400.0, 17370000.0, 17373600.0, 17377200.0, 17380800.0, 17384400.0, 17388000.0, 17391600.0, 17395200.0, 17398800.0, 17402400.0, 17406000.0, 17409600.0, 17413200.0, 17416800.0, 17420400.0, 17424000.0, 17427600.0, 17431200.0, 17434800.0, 17438400.0, 17442000.0, 17445600.0, 17449200.0, 17452800.0, 17456400.0, 17460000.0, 17463600.0, 17467200.0, 17470800.0, 17474400.0, 17478000.0, 17481600.0, 17485200.0, 17488800.0, 17492400.0, 17496000.0, 17499600.0, 17503200.0, 17506800.0, 17510400.0, 17514000.0, 17517600.0, 17521200.0, 17524800.0, 17528400.0, 17532000.0, 17535600.0, 17539200.0, 17542800.0, 17546400.0, 17550000.0, 17553600.0, 17557200.0, 17560800.0, 17564400.0, 17568000.0, 17571600.0, 17575200.0, 17578800.0, 17582400.0, 17586000.0, 17589600.0, 17593200.0, 17596800.0, 17600400.0, 17604000.0, 17607600.0, 17611200.0, 17614800.0, 17618400.0, 17622000.0, 17625600.0, 17629200.0, 17632800.0, 17636400.0, 17640000.0, 17643600.0, 17647200.0, 17650800.0, 17654400.0, 17658000.0, 17661600.0, 17665200.0, 17668800.0, 17672400.0, 17676000.0, 17679600.0, 17683200.0, 17686800.0, 17690400.0, 17694000.0, 17697600.0, 17701200.0, 17704800.0, 17708400.0, 17712000.0, 17715600.0, 17719200.0, 17722800.0, 17726400.0, 17730000.0, 17733600.0, 17737200.0, 17740800.0, 17744400.0, 17748000.0, 17751600.0, 17755200.0, 17758800.0, 17762400.0, 17766000.0, 17769600.0, 17773200.0, 17776800.0, 17780400.0, 17784000.0, 17787600.0, 17791200.0, 17794800.0, 17798400.0, 17802000.0, 17805600.0, 17809200.0, 17812800.0, 17816400.0, 17820000.0, 17823600.0, 17827200.0, 17830800.0, 17834400.0, 17838000.0, 17841600.0, 17845200.0, 17848800.0, 17852400.0, 17856000.0, 17859600.0, 17863200.0, 17866800.0, 17870400.0, 17874000.0, 17877600.0, 17881200.0, 17884800.0, 17888400.0, 17892000.0, 17895600.0, 17899200.0, 17902800.0, 17906400.0, 17910000.0, 17913600.0, 17917200.0, 17920800.0, 17924400.0, 17928000.0, 17931600.0, 17935200.0, 17938800.0, 17942400.0, 17946000.0, 17949600.0, 17953200.0, 17956800.0, 17960400.0, 17964000.0, 17967600.0, 17971200.0, 17974800.0, 17978400.0, 17982000.0, 17985600.0, 17989200.0, 17992800.0, 17996400.0, 18000000.0, 18003600.0, 18007200.0, 18010800.0, 18014400.0, 18018000.0, 18021600.0, 18025200.0, 18028800.0, 18032400.0, 18036000.0, 18039600.0, 18043200.0, 18046800.0, 18050400.0, 18054000.0, 18057600.0, 18061200.0, 18064800.0, 18068400.0, 18072000.0, 18075600.0, 18079200.0, 18082800.0, 18086400.0, 18090000.0, 18093600.0, 18097200.0, 18100800.0, 18104400.0, 18108000.0, 18111600.0, 18115200.0, 18118800.0, 18122400.0, 18126000.0, 18129600.0, 18133200.0, 18136800.0, 18140400.0, 18144000.0, 18147600.0, 18151200.0, 18154800.0, 18158400.0, 18162000.0, 18165600.0, 18169200.0, 18172800.0, 18176400.0, 18180000.0, 18183600.0, 18187200.0, 18190800.0, 18194400.0, 18198000.0, 18201600.0, 18205200.0, 18208800.0, 18212400.0, 18216000.0, 18219600.0, 18223200.0, 18226800.0, 18230400.0, 18234000.0, 18237600.0, 18241200.0, 18244800.0, 18248400.0, 18252000.0, 18255600.0, 18259200.0, 18262800.0, 18266400.0, 18270000.0, 18273600.0, 18277200.0, 18280800.0, 18284400.0, 18288000.0, 18291600.0, 18295200.0, 18298800.0, 18302400.0, 18306000.0, 18309600.0, 18313200.0, 18316800.0, 18320400.0, 18324000.0, 18327600.0, 18331200.0, 18334800.0, 18338400.0, 18342000.0, 18345600.0, 18349200.0, 18352800.0, 18356400.0, 18360000.0, 18363600.0, 18367200.0, 18370800.0, 18374400.0, 18378000.0, 18381600.0, 18385200.0, 18388800.0, 18392400.0, 18396000.0, 18399600.0, 18403200.0, 18406800.0, 18410400.0, 18414000.0, 18417600.0, 18421200.0, 18424800.0, 18428400.0, 18432000.0, 18435600.0, 18439200.0, 18442800.0, 18446400.0, 18450000.0, 18453600.0, 18457200.0, 18460800.0, 18464400.0, 18468000.0, 18471600.0, 18475200.0, 18478800.0, 18482400.0, 18486000.0, 18489600.0, 18493200.0, 18496800.0, 18500400.0, 18504000.0, 18507600.0, 18511200.0, 18514800.0, 18518400.0, 18522000.0, 18525600.0, 18529200.0, 18532800.0, 18536400.0, 18540000.0, 18543600.0, 18547200.0, 18550800.0, 18554400.0, 18558000.0, 18561600.0, 18565200.0, 18568800.0, 18572400.0, 18576000.0, 18579600.0, 18583200.0, 18586800.0, 18590400.0, 18594000.0, 18597600.0, 18601200.0, 18604800.0, 18608400.0, 18612000.0, 18615600.0, 18619200.0, 18622800.0, 18626400.0, 18630000.0, 18633600.0, 18637200.0, 18640800.0, 18644400.0, 18648000.0, 18651600.0, 18655200.0, 18658800.0, 18662400.0, 18666000.0, 18669600.0, 18673200.0, 18676800.0, 18680400.0, 18684000.0, 18687600.0, 18691200.0, 18694800.0, 18698400.0, 18702000.0, 18705600.0, 18709200.0, 18712800.0, 18716400.0, 18720000.0, 18723600.0, 18727200.0, 18730800.0, 18734400.0, 18738000.0, 18741600.0, 18745200.0, 18748800.0, 18752400.0, 18756000.0, 18759600.0, 18763200.0, 18766800.0, 18770400.0, 18774000.0, 18777600.0, 18781200.0, 18784800.0, 18788400.0, 18792000.0, 18795600.0, 18799200.0, 18802800.0, 18806400.0, 18810000.0, 18813600.0, 18817200.0, 18820800.0, 18824400.0, 18828000.0, 18831600.0, 18835200.0, 18838800.0, 18842400.0, 18846000.0, 18849600.0, 18853200.0, 18856800.0, 18860400.0, 18864000.0, 18867600.0, 18871200.0, 18874800.0, 18878400.0, 18882000.0, 18885600.0, 18889200.0, 18892800.0, 18896400.0, 18900000.0, 18903600.0, 18907200.0, 18910800.0, 18914400.0, 18918000.0, 18921600.0, 18925200.0, 18928800.0, 18932400.0, 18936000.0, 18939600.0, 18943200.0, 18946800.0, 18950400.0, 18954000.0, 18957600.0, 18961200.0, 18964800.0, 18968400.0, 18972000.0, 18975600.0, 18979200.0, 18982800.0, 18986400.0, 18990000.0, 18993600.0, 18997200.0, 19000800.0, 19004400.0, 19008000.0, 19011600.0, 19015200.0, 19018800.0, 19022400.0, 19026000.0, 19029600.0, 19033200.0, 19036800.0, 19040400.0, 19044000.0, 19047600.0, 19051200.0, 19054800.0, 19058400.0, 19062000.0, 19065600.0, 19069200.0, 19072800.0, 19076400.0, 19080000.0, 19083600.0, 19087200.0, 19090800.0, 19094400.0, 19098000.0, 19101600.0, 19105200.0, 19108800.0, 19112400.0, 19116000.0, 19119600.0, 19123200.0, 19126800.0, 19130400.0, 19134000.0, 19137600.0, 19141200.0, 19144800.0, 19148400.0, 19152000.0, 19155600.0, 19159200.0, 19162800.0, 19166400.0, 19170000.0, 19173600.0, 19177200.0, 19180800.0, 19184400.0, 19188000.0, 19191600.0, 19195200.0, 19198800.0, 19202400.0, 19206000.0, 19209600.0, 19213200.0, 19216800.0, 19220400.0, 19224000.0, 19227600.0, 19231200.0, 19234800.0, 19238400.0, 19242000.0, 19245600.0, 19249200.0, 19252800.0, 19256400.0, 19260000.0, 19263600.0, 19267200.0, 19270800.0, 19274400.0, 19278000.0, 19281600.0, 19285200.0, 19288800.0, 19292400.0, 19296000.0, 19299600.0, 19303200.0, 19306800.0, 19310400.0, 19314000.0, 19317600.0, 19321200.0, 19324800.0, 19328400.0, 19332000.0, 19335600.0, 19339200.0, 19342800.0, 19346400.0, 19350000.0, 19353600.0, 19357200.0, 19360800.0, 19364400.0, 19368000.0, 19371600.0, 19375200.0, 19378800.0, 19382400.0, 19386000.0, 19389600.0, 19393200.0, 19396800.0, 19400400.0, 19404000.0, 19407600.0, 19411200.0, 19414800.0, 19418400.0, 19422000.0, 19425600.0, 19429200.0, 19432800.0, 19436400.0, 19440000.0, 19443600.0, 19447200.0, 19450800.0, 19454400.0, 19458000.0, 19461600.0, 19465200.0, 19468800.0, 19472400.0, 19476000.0, 19479600.0, 19483200.0, 19486800.0, 19490400.0, 19494000.0, 19497600.0, 19501200.0, 19504800.0, 19508400.0, 19512000.0, 19515600.0, 19519200.0, 19522800.0, 19526400.0, 19530000.0, 19533600.0, 19537200.0, 19540800.0, 19544400.0, 19548000.0, 19551600.0, 19555200.0, 19558800.0, 19562400.0, 19566000.0, 19569600.0, 19573200.0, 19576800.0, 19580400.0, 19584000.0, 19587600.0, 19591200.0, 19594800.0, 19598400.0, 19602000.0, 19605600.0, 19609200.0, 19612800.0, 19616400.0, 19620000.0, 19623600.0, 19627200.0, 19630800.0, 19634400.0, 19638000.0, 19641600.0, 19645200.0, 19648800.0, 19652400.0, 19656000.0, 19659600.0, 19663200.0, 19666800.0, 19670400.0, 19674000.0, 19677600.0, 19681200.0, 19684800.0, 19688400.0, 19692000.0, 19695600.0, 19699200.0, 19702800.0, 19706400.0, 19710000.0, 19713600.0, 19717200.0, 19720800.0, 19724400.0, 19728000.0, 19731600.0, 19735200.0, 19738800.0, 19742400.0, 19746000.0, 19749600.0, 19753200.0, 19756800.0, 19760400.0, 19764000.0, 19767600.0, 19771200.0, 19774800.0, 19778400.0, 19782000.0, 19785600.0, 19789200.0, 19792800.0, 19796400.0, 19800000.0, 19803600.0, 19807200.0, 19810800.0, 19814400.0, 19818000.0, 19821600.0, 19825200.0, 19828800.0, 19832400.0, 19836000.0, 19839600.0, 19843200.0, 19846800.0, 19850400.0, 19854000.0, 19857600.0, 19861200.0, 19864800.0, 19868400.0, 19872000.0, 19875600.0, 19879200.0, 19882800.0, 19886400.0, 19890000.0, 19893600.0, 19897200.0, 19900800.0, 19904400.0, 19908000.0, 19911600.0, 19915200.0, 19918800.0, 19922400.0, 19926000.0, 19929600.0, 19933200.0, 19936800.0, 19940400.0, 19944000.0, 19947600.0, 19951200.0, 19954800.0, 19958400.0, 19962000.0, 19965600.0, 19969200.0, 19972800.0, 19976400.0, 19980000.0, 19983600.0, 19987200.0, 19990800.0, 19994400.0, 19998000.0, 20001600.0, 20005200.0, 20008800.0, 20012400.0, 20016000.0, 20019600.0, 20023200.0, 20026800.0, 20030400.0, 20034000.0, 20037600.0, 20041200.0, 20044800.0, 20048400.0, 20052000.0, 20055600.0, 20059200.0, 20062800.0, 20066400.0, 20070000.0, 20073600.0, 20077200.0, 20080800.0, 20084400.0, 20088000.0, 20091600.0, 20095200.0, 20098800.0, 20102400.0, 20106000.0, 20109600.0, 20113200.0, 20116800.0, 20120400.0, 20124000.0, 20127600.0, 20131200.0, 20134800.0, 20138400.0, 20142000.0, 20145600.0, 20149200.0, 20152800.0, 20156400.0, 20160000.0, 20163600.0, 20167200.0, 20170800.0, 20174400.0, 20178000.0, 20181600.0, 20185200.0, 20188800.0, 20192400.0, 20196000.0, 20199600.0, 20203200.0, 20206800.0, 20210400.0, 20214000.0, 20217600.0, 20221200.0, 20224800.0, 20228400.0, 20232000.0, 20235600.0, 20239200.0, 20242800.0, 20246400.0, 20250000.0, 20253600.0, 20257200.0, 20260800.0, 20264400.0, 20268000.0, 20271600.0, 20275200.0, 20278800.0, 20282400.0, 20286000.0, 20289600.0, 20293200.0, 20296800.0, 20300400.0, 20304000.0, 20307600.0, 20311200.0, 20314800.0, 20318400.0, 20322000.0, 20325600.0, 20329200.0, 20332800.0, 20336400.0, 20340000.0, 20343600.0, 20347200.0, 20350800.0, 20354400.0, 20358000.0, 20361600.0, 20365200.0, 20368800.0, 20372400.0, 20376000.0, 20379600.0, 20383200.0, 20386800.0, 20390400.0, 20394000.0, 20397600.0, 20401200.0, 20404800.0, 20408400.0, 20412000.0, 20415600.0, 20419200.0, 20422800.0, 20426400.0, 20430000.0, 20433600.0, 20437200.0, 20440800.0, 20444400.0, 20448000.0, 20451600.0, 20455200.0, 20458800.0, 20462400.0, 20466000.0, 20469600.0, 20473200.0, 20476800.0, 20480400.0, 20484000.0, 20487600.0, 20491200.0, 20494800.0, 20498400.0, 20502000.0, 20505600.0, 20509200.0, 20512800.0, 20516400.0, 20520000.0, 20523600.0, 20527200.0, 20530800.0, 20534400.0, 20538000.0, 20541600.0, 20545200.0, 20548800.0, 20552400.0, 20556000.0, 20559600.0, 20563200.0, 20566800.0, 20570400.0, 20574000.0, 20577600.0, 20581200.0, 20584800.0, 20588400.0, 20592000.0, 20595600.0, 20599200.0, 20602800.0, 20606400.0, 20610000.0, 20613600.0, 20617200.0, 20620800.0, 20624400.0, 20628000.0, 20631600.0, 20635200.0, 20638800.0, 20642400.0, 20646000.0, 20649600.0, 20653200.0, 20656800.0, 20660400.0, 20664000.0, 20667600.0, 20671200.0, 20674800.0, 20678400.0, 20682000.0, 20685600.0, 20689200.0, 20692800.0, 20696400.0, 20700000.0, 20703600.0, 20707200.0, 20710800.0, 20714400.0, 20718000.0, 20721600.0, 20725200.0, 20728800.0, 20732400.0, 20736000.0, 20739600.0, 20743200.0, 20746800.0, 20750400.0, 20754000.0, 20757600.0, 20761200.0, 20764800.0, 20768400.0, 20772000.0, 20775600.0, 20779200.0, 20782800.0, 20786400.0, 20790000.0, 20793600.0, 20797200.0, 20800800.0, 20804400.0, 20808000.0, 20811600.0, 20815200.0, 20818800.0, 20822400.0, 20826000.0, 20829600.0, 20833200.0, 20836800.0, 20840400.0, 20844000.0, 20847600.0, 20851200.0, 20854800.0, 20858400.0, 20862000.0, 20865600.0, 20869200.0, 20872800.0, 20876400.0, 20880000.0, 20883600.0, 20887200.0, 20890800.0, 20894400.0, 20898000.0, 20901600.0, 20905200.0, 20908800.0, 20912400.0, 20916000.0, 20919600.0, 20923200.0, 20926800.0, 20930400.0, 20934000.0, 20937600.0, 20941200.0, 20944800.0, 20948400.0, 20952000.0, 20955600.0, 20959200.0, 20962800.0, 20966400.0, 20970000.0, 20973600.0, 20977200.0, 20980800.0, 20984400.0, 20988000.0, 20991600.0, 20995200.0, 20998800.0, 21002400.0, 21006000.0, 21009600.0, 21013200.0, 21016800.0, 21020400.0, 21024000.0, 21027600.0, 21031200.0, 21034800.0, 21038400.0, 21042000.0, 21045600.0, 21049200.0, 21052800.0, 21056400.0, 21060000.0, 21063600.0, 21067200.0, 21070800.0, 21074400.0, 21078000.0, 21081600.0, 21085200.0, 21088800.0, 21092400.0, 21096000.0, 21099600.0, 21103200.0, 21106800.0, 21110400.0, 21114000.0, 21117600.0, 21121200.0, 21124800.0, 21128400.0, 21132000.0, 21135600.0, 21139200.0, 21142800.0, 21146400.0, 21150000.0, 21153600.0, 21157200.0, 21160800.0, 21164400.0, 21168000.0, 21171600.0, 21175200.0, 21178800.0, 21182400.0, 21186000.0, 21189600.0, 21193200.0, 21196800.0, 21200400.0, 21204000.0, 21207600.0, 21211200.0, 21214800.0, 21218400.0, 21222000.0, 21225600.0, 21229200.0, 21232800.0, 21236400.0, 21240000.0, 21243600.0, 21247200.0, 21250800.0, 21254400.0, 21258000.0, 21261600.0, 21265200.0, 21268800.0, 21272400.0, 21276000.0, 21279600.0, 21283200.0, 21286800.0, 21290400.0, 21294000.0, 21297600.0, 21301200.0, 21304800.0, 21308400.0, 21312000.0, 21315600.0, 21319200.0, 21322800.0, 21326400.0, 21330000.0, 21333600.0, 21337200.0, 21340800.0, 21344400.0, 21348000.0, 21351600.0, 21355200.0, 21358800.0, 21362400.0, 21366000.0, 21369600.0, 21373200.0, 21376800.0, 21380400.0, 21384000.0, 21387600.0, 21391200.0, 21394800.0, 21398400.0, 21402000.0, 21405600.0, 21409200.0, 21412800.0, 21416400.0, 21420000.0, 21423600.0, 21427200.0, 21430800.0, 21434400.0, 21438000.0, 21441600.0, 21445200.0, 21448800.0, 21452400.0, 21456000.0, 21459600.0, 21463200.0, 21466800.0, 21470400.0, 21474000.0, 21477600.0, 21481200.0, 21484800.0, 21488400.0, 21492000.0, 21495600.0, 21499200.0, 21502800.0, 21506400.0, 21510000.0, 21513600.0, 21517200.0, 21520800.0, 21524400.0, 21528000.0, 21531600.0, 21535200.0, 21538800.0, 21542400.0, 21546000.0, 21549600.0, 21553200.0, 21556800.0, 21560400.0, 21564000.0, 21567600.0, 21571200.0, 21574800.0, 21578400.0, 21582000.0, 21585600.0, 21589200.0, 21592800.0, 21596400.0, 21600000.0, 21603600.0, 21607200.0, 21610800.0, 21614400.0, 21618000.0, 21621600.0, 21625200.0, 21628800.0, 21632400.0, 21636000.0, 21639600.0, 21643200.0, 21646800.0, 21650400.0, 21654000.0, 21657600.0, 21661200.0, 21664800.0, 21668400.0, 21672000.0, 21675600.0, 21679200.0, 21682800.0, 21686400.0, 21690000.0, 21693600.0, 21697200.0, 21700800.0, 21704400.0, 21708000.0, 21711600.0, 21715200.0, 21718800.0, 21722400.0, 21726000.0, 21729600.0, 21733200.0, 21736800.0, 21740400.0, 21744000.0, 21747600.0, 21751200.0, 21754800.0, 21758400.0, 21762000.0, 21765600.0, 21769200.0, 21772800.0, 21776400.0, 21780000.0, 21783600.0, 21787200.0, 21790800.0, 21794400.0, 21798000.0, 21801600.0, 21805200.0, 21808800.0, 21812400.0, 21816000.0, 21819600.0, 21823200.0, 21826800.0, 21830400.0, 21834000.0, 21837600.0, 21841200.0, 21844800.0, 21848400.0, 21852000.0, 21855600.0, 21859200.0, 21862800.0, 21866400.0, 21870000.0, 21873600.0, 21877200.0, 21880800.0, 21884400.0, 21888000.0, 21891600.0, 21895200.0, 21898800.0, 21902400.0, 21906000.0, 21909600.0, 21913200.0, 21916800.0, 21920400.0, 21924000.0, 21927600.0, 21931200.0, 21934800.0, 21938400.0, 21942000.0, 21945600.0, 21949200.0, 21952800.0, 21956400.0, 21960000.0, 21963600.0, 21967200.0, 21970800.0, 21974400.0, 21978000.0, 21981600.0, 21985200.0, 21988800.0, 21992400.0, 21996000.0, 21999600.0, 22003200.0, 22006800.0, 22010400.0, 22014000.0, 22017600.0, 22021200.0, 22024800.0, 22028400.0, 22032000.0, 22035600.0, 22039200.0, 22042800.0, 22046400.0, 22050000.0, 22053600.0, 22057200.0, 22060800.0, 22064400.0, 22068000.0, 22071600.0, 22075200.0, 22078800.0, 22082400.0, 22086000.0, 22089600.0, 22093200.0, 22096800.0, 22100400.0, 22104000.0, 22107600.0, 22111200.0, 22114800.0, 22118400.0, 22122000.0, 22125600.0, 22129200.0, 22132800.0, 22136400.0, 22140000.0, 22143600.0, 22147200.0, 22150800.0, 22154400.0, 22158000.0, 22161600.0, 22165200.0, 22168800.0, 22172400.0, 22176000.0, 22179600.0, 22183200.0, 22186800.0, 22190400.0, 22194000.0, 22197600.0, 22201200.0, 22204800.0, 22208400.0, 22212000.0, 22215600.0, 22219200.0, 22222800.0, 22226400.0, 22230000.0, 22233600.0, 22237200.0, 22240800.0, 22244400.0, 22248000.0, 22251600.0, 22255200.0, 22258800.0, 22262400.0, 22266000.0, 22269600.0, 22273200.0, 22276800.0, 22280400.0, 22284000.0, 22287600.0, 22291200.0, 22294800.0, 22298400.0, 22302000.0, 22305600.0, 22309200.0, 22312800.0, 22316400.0, 22320000.0, 22323600.0, 22327200.0, 22330800.0, 22334400.0, 22338000.0, 22341600.0, 22345200.0, 22348800.0, 22352400.0, 22356000.0, 22359600.0, 22363200.0, 22366800.0, 22370400.0, 22374000.0, 22377600.0, 22381200.0, 22384800.0, 22388400.0, 22392000.0, 22395600.0, 22399200.0, 22402800.0, 22406400.0, 22410000.0, 22413600.0, 22417200.0, 22420800.0, 22424400.0, 22428000.0, 22431600.0, 22435200.0, 22438800.0, 22442400.0, 22446000.0, 22449600.0, 22453200.0, 22456800.0, 22460400.0, 22464000.0, 22467600.0, 22471200.0, 22474800.0, 22478400.0, 22482000.0, 22485600.0, 22489200.0, 22492800.0, 22496400.0, 22500000.0, 22503600.0, 22507200.0, 22510800.0, 22514400.0, 22518000.0, 22521600.0, 22525200.0, 22528800.0, 22532400.0, 22536000.0, 22539600.0, 22543200.0, 22546800.0, 22550400.0, 22554000.0, 22557600.0, 22561200.0, 22564800.0, 22568400.0, 22572000.0, 22575600.0, 22579200.0, 22582800.0, 22586400.0, 22590000.0, 22593600.0, 22597200.0, 22600800.0, 22604400.0, 22608000.0, 22611600.0, 22615200.0, 22618800.0, 22622400.0, 22626000.0, 22629600.0, 22633200.0, 22636800.0, 22640400.0, 22644000.0, 22647600.0, 22651200.0, 22654800.0, 22658400.0, 22662000.0, 22665600.0, 22669200.0, 22672800.0, 22676400.0, 22680000.0, 22683600.0, 22687200.0, 22690800.0, 22694400.0, 22698000.0, 22701600.0, 22705200.0, 22708800.0, 22712400.0, 22716000.0, 22719600.0, 22723200.0, 22726800.0, 22730400.0, 22734000.0, 22737600.0, 22741200.0, 22744800.0, 22748400.0, 22752000.0, 22755600.0, 22759200.0, 22762800.0, 22766400.0, 22770000.0, 22773600.0, 22777200.0, 22780800.0, 22784400.0, 22788000.0, 22791600.0, 22795200.0, 22798800.0, 22802400.0, 22806000.0, 22809600.0, 22813200.0, 22816800.0, 22820400.0, 22824000.0, 22827600.0, 22831200.0, 22834800.0, 22838400.0, 22842000.0, 22845600.0, 22849200.0, 22852800.0, 22856400.0, 22860000.0, 22863600.0, 22867200.0, 22870800.0, 22874400.0, 22878000.0, 22881600.0, 22885200.0, 22888800.0, 22892400.0, 22896000.0, 22899600.0, 22903200.0, 22906800.0, 22910400.0, 22914000.0, 22917600.0, 22921200.0, 22924800.0, 22928400.0, 22932000.0, 22935600.0, 22939200.0, 22942800.0, 22946400.0, 22950000.0, 22953600.0, 22957200.0, 22960800.0, 22964400.0, 22968000.0, 22971600.0, 22975200.0, 22978800.0, 22982400.0, 22986000.0, 22989600.0, 22993200.0, 22996800.0, 23000400.0, 23004000.0, 23007600.0, 23011200.0, 23014800.0, 23018400.0, 23022000.0, 23025600.0, 23029200.0, 23032800.0, 23036400.0, 23040000.0, 23043600.0, 23047200.0, 23050800.0, 23054400.0, 23058000.0, 23061600.0, 23065200.0, 23068800.0, 23072400.0, 23076000.0, 23079600.0, 23083200.0, 23086800.0, 23090400.0, 23094000.0, 23097600.0, 23101200.0, 23104800.0, 23108400.0, 23112000.0, 23115600.0, 23119200.0, 23122800.0, 23126400.0, 23130000.0, 23133600.0, 23137200.0, 23140800.0, 23144400.0, 23148000.0, 23151600.0, 23155200.0, 23158800.0, 23162400.0, 23166000.0, 23169600.0, 23173200.0, 23176800.0, 23180400.0, 23184000.0, 23187600.0, 23191200.0, 23194800.0, 23198400.0, 23202000.0, 23205600.0, 23209200.0, 23212800.0, 23216400.0, 23220000.0, 23223600.0, 23227200.0, 23230800.0, 23234400.0, 23238000.0, 23241600.0, 23245200.0, 23248800.0, 23252400.0, 23256000.0, 23259600.0, 23263200.0, 23266800.0, 23270400.0, 23274000.0, 23277600.0, 23281200.0, 23284800.0, 23288400.0, 23292000.0, 23295600.0, 23299200.0, 23302800.0, 23306400.0, 23310000.0, 23313600.0, 23317200.0, 23320800.0, 23324400.0, 23328000.0, 23331600.0, 23335200.0, 23338800.0, 23342400.0, 23346000.0, 23349600.0, 23353200.0, 23356800.0, 23360400.0, 23364000.0, 23367600.0, 23371200.0, 23374800.0, 23378400.0, 23382000.0, 23385600.0, 23389200.0, 23392800.0, 23396400.0, 23400000.0, 23403600.0, 23407200.0, 23410800.0, 23414400.0, 23418000.0, 23421600.0, 23425200.0, 23428800.0, 23432400.0, 23436000.0, 23439600.0, 23443200.0, 23446800.0, 23450400.0, 23454000.0, 23457600.0, 23461200.0, 23464800.0, 23468400.0, 23472000.0, 23475600.0, 23479200.0, 23482800.0, 23486400.0, 23490000.0, 23493600.0, 23497200.0, 23500800.0, 23504400.0, 23508000.0, 23511600.0, 23515200.0, 23518800.0, 23522400.0, 23526000.0, 23529600.0, 23533200.0, 23536800.0, 23540400.0, 23544000.0, 23547600.0, 23551200.0, 23554800.0, 23558400.0, 23562000.0, 23565600.0, 23569200.0, 23572800.0, 23576400.0, 23580000.0, 23583600.0, 23587200.0, 23590800.0, 23594400.0, 23598000.0, 23601600.0, 23605200.0, 23608800.0, 23612400.0, 23616000.0, 23619600.0, 23623200.0, 23626800.0, 23630400.0, 23634000.0, 23637600.0, 23641200.0, 23644800.0, 23648400.0, 23652000.0, 23655600.0, 23659200.0, 23662800.0, 23666400.0, 23670000.0, 23673600.0, 23677200.0, 23680800.0, 23684400.0, 23688000.0, 23691600.0, 23695200.0, 23698800.0, 23702400.0, 23706000.0, 23709600.0, 23713200.0, 23716800.0, 23720400.0, 23724000.0, 23727600.0, 23731200.0, 23734800.0, 23738400.0, 23742000.0, 23745600.0, 23749200.0, 23752800.0, 23756400.0, 23760000.0, 23763600.0, 23767200.0, 23770800.0, 23774400.0, 23778000.0, 23781600.0, 23785200.0, 23788800.0, 23792400.0, 23796000.0, 23799600.0, 23803200.0, 23806800.0, 23810400.0, 23814000.0, 23817600.0, 23821200.0, 23824800.0, 23828400.0, 23832000.0, 23835600.0, 23839200.0, 23842800.0, 23846400.0, 23850000.0, 23853600.0, 23857200.0, 23860800.0, 23864400.0, 23868000.0, 23871600.0, 23875200.0, 23878800.0, 23882400.0, 23886000.0, 23889600.0, 23893200.0, 23896800.0, 23900400.0, 23904000.0, 23907600.0, 23911200.0, 23914800.0, 23918400.0, 23922000.0, 23925600.0, 23929200.0, 23932800.0, 23936400.0, 23940000.0, 23943600.0, 23947200.0, 23950800.0, 23954400.0, 23958000.0, 23961600.0, 23965200.0, 23968800.0, 23972400.0, 23976000.0, 23979600.0, 23983200.0, 23986800.0, 23990400.0, 23994000.0, 23997600.0, 24001200.0, 24004800.0, 24008400.0, 24012000.0, 24015600.0, 24019200.0, 24022800.0, 24026400.0, 24030000.0, 24033600.0, 24037200.0, 24040800.0, 24044400.0, 24048000.0, 24051600.0, 24055200.0, 24058800.0, 24062400.0, 24066000.0, 24069600.0, 24073200.0, 24076800.0, 24080400.0, 24084000.0, 24087600.0, 24091200.0, 24094800.0, 24098400.0, 24102000.0, 24105600.0, 24109200.0, 24112800.0, 24116400.0, 24120000.0, 24123600.0, 24127200.0, 24130800.0, 24134400.0, 24138000.0, 24141600.0, 24145200.0, 24148800.0, 24152400.0, 24156000.0, 24159600.0, 24163200.0, 24166800.0, 24170400.0, 24174000.0, 24177600.0, 24181200.0, 24184800.0, 24188400.0, 24192000.0, 24195600.0, 24199200.0, 24202800.0, 24206400.0, 24210000.0, 24213600.0, 24217200.0, 24220800.0, 24224400.0, 24228000.0, 24231600.0, 24235200.0, 24238800.0, 24242400.0, 24246000.0, 24249600.0, 24253200.0, 24256800.0, 24260400.0, 24264000.0, 24267600.0, 24271200.0, 24274800.0, 24278400.0, 24282000.0, 24285600.0, 24289200.0, 24292800.0, 24296400.0, 24300000.0, 24303600.0, 24307200.0, 24310800.0, 24314400.0, 24318000.0, 24321600.0, 24325200.0, 24328800.0, 24332400.0, 24336000.0, 24339600.0, 24343200.0, 24346800.0, 24350400.0, 24354000.0, 24357600.0, 24361200.0, 24364800.0, 24368400.0, 24372000.0, 24375600.0, 24379200.0, 24382800.0, 24386400.0, 24390000.0, 24393600.0, 24397200.0, 24400800.0, 24404400.0, 24408000.0, 24411600.0, 24415200.0, 24418800.0, 24422400.0, 24426000.0, 24429600.0, 24433200.0, 24436800.0, 24440400.0, 24444000.0, 24447600.0, 24451200.0, 24454800.0, 24458400.0, 24462000.0, 24465600.0, 24469200.0, 24472800.0, 24476400.0, 24480000.0, 24483600.0, 24487200.0, 24490800.0, 24494400.0, 24498000.0, 24501600.0, 24505200.0, 24508800.0, 24512400.0, 24516000.0, 24519600.0, 24523200.0, 24526800.0, 24530400.0, 24534000.0, 24537600.0, 24541200.0, 24544800.0, 24548400.0, 24552000.0, 24555600.0, 24559200.0, 24562800.0, 24566400.0, 24570000.0, 24573600.0, 24577200.0, 24580800.0, 24584400.0, 24588000.0, 24591600.0, 24595200.0, 24598800.0, 24602400.0, 24606000.0, 24609600.0, 24613200.0, 24616800.0, 24620400.0, 24624000.0, 24627600.0, 24631200.0, 24634800.0, 24638400.0, 24642000.0, 24645600.0, 24649200.0, 24652800.0, 24656400.0, 24660000.0, 24663600.0, 24667200.0, 24670800.0, 24674400.0, 24678000.0, 24681600.0, 24685200.0, 24688800.0, 24692400.0, 24696000.0, 24699600.0, 24703200.0, 24706800.0, 24710400.0, 24714000.0, 24717600.0, 24721200.0, 24724800.0, 24728400.0, 24732000.0, 24735600.0, 24739200.0, 24742800.0, 24746400.0, 24750000.0, 24753600.0, 24757200.0, 24760800.0, 24764400.0, 24768000.0, 24771600.0, 24775200.0, 24778800.0, 24782400.0, 24786000.0, 24789600.0, 24793200.0, 24796800.0, 24800400.0, 24804000.0, 24807600.0, 24811200.0, 24814800.0, 24818400.0, 24822000.0, 24825600.0, 24829200.0, 24832800.0, 24836400.0, 24840000.0, 24843600.0, 24847200.0, 24850800.0, 24854400.0, 24858000.0, 24861600.0, 24865200.0, 24868800.0, 24872400.0, 24876000.0, 24879600.0, 24883200.0, 24886800.0, 24890400.0, 24894000.0, 24897600.0, 24901200.0, 24904800.0, 24908400.0, 24912000.0, 24915600.0, 24919200.0, 24922800.0, 24926400.0, 24930000.0, 24933600.0, 24937200.0, 24940800.0, 24944400.0, 24948000.0, 24951600.0, 24955200.0, 24958800.0, 24962400.0, 24966000.0, 24969600.0, 24973200.0, 24976800.0, 24980400.0, 24984000.0, 24987600.0, 24991200.0, 24994800.0, 24998400.0, 25002000.0, 25005600.0, 25009200.0, 25012800.0, 25016400.0, 25020000.0, 25023600.0, 25027200.0, 25030800.0, 25034400.0, 25038000.0, 25041600.0, 25045200.0, 25048800.0, 25052400.0, 25056000.0, 25059600.0, 25063200.0, 25066800.0, 25070400.0, 25074000.0, 25077600.0, 25081200.0, 25084800.0, 25088400.0, 25092000.0, 25095600.0, 25099200.0, 25102800.0, 25106400.0, 25110000.0, 25113600.0, 25117200.0, 25120800.0, 25124400.0, 25128000.0, 25131600.0, 25135200.0, 25138800.0, 25142400.0, 25146000.0, 25149600.0, 25153200.0, 25156800.0, 25160400.0, 25164000.0, 25167600.0, 25171200.0, 25174800.0, 25178400.0, 25182000.0, 25185600.0, 25189200.0, 25192800.0, 25196400.0, 25200000.0, 25203600.0, 25207200.0, 25210800.0, 25214400.0, 25218000.0, 25221600.0, 25225200.0, 25228800.0, 25232400.0, 25236000.0, 25239600.0, 25243200.0, 25246800.0, 25250400.0, 25254000.0, 25257600.0, 25261200.0, 25264800.0, 25268400.0, 25272000.0, 25275600.0, 25279200.0, 25282800.0, 25286400.0, 25290000.0, 25293600.0, 25297200.0, 25300800.0, 25304400.0, 25308000.0, 25311600.0, 25315200.0, 25318800.0, 25322400.0, 25326000.0, 25329600.0, 25333200.0, 25336800.0, 25340400.0, 25344000.0, 25347600.0, 25351200.0, 25354800.0, 25358400.0, 25362000.0, 25365600.0, 25369200.0, 25372800.0, 25376400.0, 25380000.0, 25383600.0, 25387200.0, 25390800.0, 25394400.0, 25398000.0, 25401600.0, 25405200.0, 25408800.0, 25412400.0, 25416000.0, 25419600.0, 25423200.0, 25426800.0, 25430400.0, 25434000.0, 25437600.0, 25441200.0, 25444800.0, 25448400.0, 25452000.0, 25455600.0, 25459200.0, 25462800.0, 25466400.0, 25470000.0, 25473600.0, 25477200.0, 25480800.0, 25484400.0, 25488000.0, 25491600.0, 25495200.0, 25498800.0, 25502400.0, 25506000.0, 25509600.0, 25513200.0, 25516800.0, 25520400.0, 25524000.0, 25527600.0, 25531200.0, 25534800.0, 25538400.0, 25542000.0, 25545600.0, 25549200.0, 25552800.0, 25556400.0, 25560000.0, 25563600.0, 25567200.0, 25570800.0, 25574400.0, 25578000.0, 25581600.0, 25585200.0, 25588800.0, 25592400.0, 25596000.0, 25599600.0, 25603200.0, 25606800.0, 25610400.0, 25614000.0, 25617600.0, 25621200.0, 25624800.0, 25628400.0, 25632000.0, 25635600.0, 25639200.0, 25642800.0, 25646400.0, 25650000.0, 25653600.0, 25657200.0, 25660800.0, 25664400.0, 25668000.0, 25671600.0, 25675200.0, 25678800.0, 25682400.0, 25686000.0, 25689600.0, 25693200.0, 25696800.0, 25700400.0, 25704000.0, 25707600.0, 25711200.0, 25714800.0, 25718400.0, 25722000.0, 25725600.0, 25729200.0, 25732800.0, 25736400.0, 25740000.0, 25743600.0, 25747200.0, 25750800.0, 25754400.0, 25758000.0, 25761600.0, 25765200.0, 25768800.0, 25772400.0, 25776000.0, 25779600.0, 25783200.0, 25786800.0, 25790400.0, 25794000.0, 25797600.0, 25801200.0, 25804800.0, 25808400.0, 25812000.0, 25815600.0, 25819200.0, 25822800.0, 25826400.0, 25830000.0, 25833600.0, 25837200.0, 25840800.0, 25844400.0, 25848000.0, 25851600.0, 25855200.0, 25858800.0, 25862400.0, 25866000.0, 25869600.0, 25873200.0, 25876800.0, 25880400.0, 25884000.0, 25887600.0, 25891200.0, 25894800.0, 25898400.0, 25902000.0, 25905600.0, 25909200.0, 25912800.0, 25916400.0, 25920000.0, 25923600.0, 25927200.0, 25930800.0, 25934400.0, 25938000.0, 25941600.0, 25945200.0, 25948800.0, 25952400.0, 25956000.0, 25959600.0, 25963200.0, 25966800.0, 25970400.0, 25974000.0, 25977600.0, 25981200.0, 25984800.0, 25988400.0, 25992000.0, 25995600.0, 25999200.0, 26002800.0, 26006400.0, 26010000.0, 26013600.0, 26017200.0, 26020800.0, 26024400.0, 26028000.0, 26031600.0, 26035200.0, 26038800.0, 26042400.0, 26046000.0, 26049600.0, 26053200.0, 26056800.0, 26060400.0, 26064000.0, 26067600.0, 26071200.0, 26074800.0, 26078400.0, 26082000.0, 26085600.0, 26089200.0, 26092800.0, 26096400.0, 26100000.0, 26103600.0, 26107200.0, 26110800.0, 26114400.0, 26118000.0, 26121600.0, 26125200.0, 26128800.0, 26132400.0, 26136000.0, 26139600.0, 26143200.0, 26146800.0, 26150400.0, 26154000.0, 26157600.0, 26161200.0, 26164800.0, 26168400.0, 26172000.0, 26175600.0, 26179200.0, 26182800.0, 26186400.0, 26190000.0, 26193600.0, 26197200.0, 26200800.0, 26204400.0, 26208000.0, 26211600.0, 26215200.0, 26218800.0, 26222400.0, 26226000.0, 26229600.0, 26233200.0, 26236800.0, 26240400.0, 26244000.0, 26247600.0, 26251200.0, 26254800.0, 26258400.0, 26262000.0, 26265600.0, 26269200.0, 26272800.0, 26276400.0, 26280000.0, 26283600.0, 26287200.0, 26290800.0, 26294400.0, 26298000.0, 26301600.0, 26305200.0, 26308800.0, 26312400.0, 26316000.0, 26319600.0, 26323200.0, 26326800.0, 26330400.0, 26334000.0, 26337600.0, 26341200.0, 26344800.0, 26348400.0, 26352000.0, 26355600.0, 26359200.0, 26362800.0, 26366400.0, 26370000.0, 26373600.0, 26377200.0, 26380800.0, 26384400.0, 26388000.0, 26391600.0, 26395200.0, 26398800.0, 26402400.0, 26406000.0, 26409600.0, 26413200.0, 26416800.0, 26420400.0, 26424000.0, 26427600.0, 26431200.0, 26434800.0, 26438400.0, 26442000.0, 26445600.0, 26449200.0, 26452800.0, 26456400.0, 26460000.0, 26463600.0, 26467200.0, 26470800.0, 26474400.0, 26478000.0, 26481600.0, 26485200.0, 26488800.0, 26492400.0, 26496000.0, 26499600.0, 26503200.0, 26506800.0, 26510400.0, 26514000.0, 26517600.0, 26521200.0, 26524800.0, 26528400.0, 26532000.0, 26535600.0, 26539200.0, 26542800.0, 26546400.0, 26550000.0, 26553600.0, 26557200.0, 26560800.0, 26564400.0, 26568000.0, 26571600.0, 26575200.0, 26578800.0, 26582400.0, 26586000.0, 26589600.0, 26593200.0, 26596800.0, 26600400.0, 26604000.0, 26607600.0, 26611200.0, 26614800.0, 26618400.0, 26622000.0, 26625600.0, 26629200.0, 26632800.0, 26636400.0, 26640000.0, 26643600.0, 26647200.0, 26650800.0, 26654400.0, 26658000.0, 26661600.0, 26665200.0, 26668800.0, 26672400.0, 26676000.0, 26679600.0, 26683200.0, 26686800.0, 26690400.0, 26694000.0, 26697600.0, 26701200.0, 26704800.0, 26708400.0, 26712000.0, 26715600.0, 26719200.0, 26722800.0, 26726400.0, 26730000.0, 26733600.0, 26737200.0, 26740800.0, 26744400.0, 26748000.0, 26751600.0, 26755200.0, 26758800.0, 26762400.0, 26766000.0, 26769600.0, 26773200.0, 26776800.0, 26780400.0, 26784000.0, 26787600.0, 26791200.0, 26794800.0, 26798400.0, 26802000.0, 26805600.0, 26809200.0, 26812800.0, 26816400.0, 26820000.0, 26823600.0, 26827200.0, 26830800.0, 26834400.0, 26838000.0, 26841600.0, 26845200.0, 26848800.0, 26852400.0, 26856000.0, 26859600.0, 26863200.0, 26866800.0, 26870400.0, 26874000.0, 26877600.0, 26881200.0, 26884800.0, 26888400.0, 26892000.0, 26895600.0, 26899200.0, 26902800.0, 26906400.0, 26910000.0, 26913600.0, 26917200.0, 26920800.0, 26924400.0, 26928000.0, 26931600.0, 26935200.0, 26938800.0, 26942400.0, 26946000.0, 26949600.0, 26953200.0, 26956800.0, 26960400.0, 26964000.0, 26967600.0, 26971200.0, 26974800.0, 26978400.0, 26982000.0, 26985600.0, 26989200.0, 26992800.0, 26996400.0, 27000000.0, 27003600.0, 27007200.0, 27010800.0, 27014400.0, 27018000.0, 27021600.0, 27025200.0, 27028800.0, 27032400.0, 27036000.0, 27039600.0, 27043200.0, 27046800.0, 27050400.0, 27054000.0, 27057600.0, 27061200.0, 27064800.0, 27068400.0, 27072000.0, 27075600.0, 27079200.0, 27082800.0, 27086400.0, 27090000.0, 27093600.0, 27097200.0, 27100800.0, 27104400.0, 27108000.0, 27111600.0, 27115200.0, 27118800.0, 27122400.0, 27126000.0, 27129600.0, 27133200.0, 27136800.0, 27140400.0, 27144000.0, 27147600.0, 27151200.0, 27154800.0, 27158400.0, 27162000.0, 27165600.0, 27169200.0, 27172800.0, 27176400.0, 27180000.0, 27183600.0, 27187200.0, 27190800.0, 27194400.0, 27198000.0, 27201600.0, 27205200.0, 27208800.0, 27212400.0, 27216000.0, 27219600.0, 27223200.0, 27226800.0, 27230400.0, 27234000.0, 27237600.0, 27241200.0, 27244800.0, 27248400.0, 27252000.0, 27255600.0, 27259200.0, 27262800.0, 27266400.0, 27270000.0, 27273600.0, 27277200.0, 27280800.0, 27284400.0, 27288000.0, 27291600.0, 27295200.0, 27298800.0, 27302400.0, 27306000.0, 27309600.0, 27313200.0, 27316800.0, 27320400.0, 27324000.0, 27327600.0, 27331200.0, 27334800.0, 27338400.0, 27342000.0, 27345600.0, 27349200.0, 27352800.0, 27356400.0, 27360000.0, 27363600.0, 27367200.0, 27370800.0, 27374400.0, 27378000.0, 27381600.0, 27385200.0, 27388800.0, 27392400.0, 27396000.0, 27399600.0, 27403200.0, 27406800.0, 27410400.0, 27414000.0, 27417600.0, 27421200.0, 27424800.0, 27428400.0, 27432000.0, 27435600.0, 27439200.0, 27442800.0, 27446400.0, 27450000.0, 27453600.0, 27457200.0, 27460800.0, 27464400.0, 27468000.0, 27471600.0, 27475200.0, 27478800.0, 27482400.0, 27486000.0, 27489600.0, 27493200.0, 27496800.0, 27500400.0, 27504000.0, 27507600.0, 27511200.0, 27514800.0, 27518400.0, 27522000.0, 27525600.0, 27529200.0, 27532800.0, 27536400.0, 27540000.0, 27543600.0, 27547200.0, 27550800.0, 27554400.0, 27558000.0, 27561600.0, 27565200.0, 27568800.0, 27572400.0, 27576000.0, 27579600.0, 27583200.0, 27586800.0, 27590400.0, 27594000.0, 27597600.0, 27601200.0, 27604800.0, 27608400.0, 27612000.0, 27615600.0, 27619200.0, 27622800.0, 27626400.0, 27630000.0, 27633600.0, 27637200.0, 27640800.0, 27644400.0, 27648000.0, 27651600.0, 27655200.0, 27658800.0, 27662400.0, 27666000.0, 27669600.0, 27673200.0, 27676800.0, 27680400.0, 27684000.0, 27687600.0, 27691200.0, 27694800.0, 27698400.0, 27702000.0, 27705600.0, 27709200.0, 27712800.0, 27716400.0, 27720000.0, 27723600.0, 27727200.0, 27730800.0, 27734400.0, 27738000.0, 27741600.0, 27745200.0, 27748800.0, 27752400.0, 27756000.0, 27759600.0, 27763200.0, 27766800.0, 27770400.0, 27774000.0, 27777600.0, 27781200.0, 27784800.0, 27788400.0, 27792000.0, 27795600.0, 27799200.0, 27802800.0, 27806400.0, 27810000.0, 27813600.0, 27817200.0, 27820800.0, 27824400.0, 27828000.0, 27831600.0, 27835200.0, 27838800.0, 27842400.0, 27846000.0, 27849600.0, 27853200.0, 27856800.0, 27860400.0, 27864000.0, 27867600.0, 27871200.0, 27874800.0, 27878400.0, 27882000.0, 27885600.0, 27889200.0, 27892800.0, 27896400.0, 27900000.0, 27903600.0, 27907200.0, 27910800.0, 27914400.0, 27918000.0, 27921600.0, 27925200.0, 27928800.0, 27932400.0, 27936000.0, 27939600.0, 27943200.0, 27946800.0, 27950400.0, 27954000.0, 27957600.0, 27961200.0, 27964800.0, 27968400.0, 27972000.0, 27975600.0, 27979200.0, 27982800.0, 27986400.0, 27990000.0, 27993600.0, 27997200.0, 28000800.0, 28004400.0, 28008000.0, 28011600.0, 28015200.0, 28018800.0, 28022400.0, 28026000.0, 28029600.0, 28033200.0, 28036800.0, 28040400.0, 28044000.0, 28047600.0, 28051200.0, 28054800.0, 28058400.0, 28062000.0, 28065600.0, 28069200.0, 28072800.0, 28076400.0, 28080000.0, 28083600.0, 28087200.0, 28090800.0, 28094400.0, 28098000.0, 28101600.0, 28105200.0, 28108800.0, 28112400.0, 28116000.0, 28119600.0, 28123200.0, 28126800.0, 28130400.0, 28134000.0, 28137600.0, 28141200.0, 28144800.0, 28148400.0, 28152000.0, 28155600.0, 28159200.0, 28162800.0, 28166400.0, 28170000.0, 28173600.0, 28177200.0, 28180800.0, 28184400.0, 28188000.0, 28191600.0, 28195200.0, 28198800.0, 28202400.0, 28206000.0, 28209600.0, 28213200.0, 28216800.0, 28220400.0, 28224000.0, 28227600.0, 28231200.0, 28234800.0, 28238400.0, 28242000.0, 28245600.0, 28249200.0, 28252800.0, 28256400.0, 28260000.0, 28263600.0, 28267200.0, 28270800.0, 28274400.0, 28278000.0, 28281600.0, 28285200.0, 28288800.0, 28292400.0, 28296000.0, 28299600.0, 28303200.0, 28306800.0, 28310400.0, 28314000.0, 28317600.0, 28321200.0, 28324800.0, 28328400.0, 28332000.0, 28335600.0, 28339200.0, 28342800.0, 28346400.0, 28350000.0, 28353600.0, 28357200.0, 28360800.0, 28364400.0, 28368000.0, 28371600.0, 28375200.0, 28378800.0, 28382400.0, 28386000.0, 28389600.0, 28393200.0, 28396800.0, 28400400.0, 28404000.0, 28407600.0, 28411200.0, 28414800.0, 28418400.0, 28422000.0, 28425600.0, 28429200.0, 28432800.0, 28436400.0, 28440000.0, 28443600.0, 28447200.0, 28450800.0, 28454400.0, 28458000.0, 28461600.0, 28465200.0, 28468800.0, 28472400.0, 28476000.0, 28479600.0, 28483200.0, 28486800.0, 28490400.0, 28494000.0, 28497600.0, 28501200.0, 28504800.0, 28508400.0, 28512000.0, 28515600.0, 28519200.0, 28522800.0, 28526400.0, 28530000.0, 28533600.0, 28537200.0, 28540800.0, 28544400.0, 28548000.0, 28551600.0, 28555200.0, 28558800.0, 28562400.0, 28566000.0, 28569600.0, 28573200.0, 28576800.0, 28580400.0, 28584000.0, 28587600.0, 28591200.0, 28594800.0, 28598400.0, 28602000.0, 28605600.0, 28609200.0, 28612800.0, 28616400.0, 28620000.0, 28623600.0, 28627200.0, 28630800.0, 28634400.0, 28638000.0, 28641600.0, 28645200.0, 28648800.0, 28652400.0, 28656000.0, 28659600.0, 28663200.0, 28666800.0, 28670400.0, 28674000.0, 28677600.0, 28681200.0, 28684800.0, 28688400.0, 28692000.0, 28695600.0, 28699200.0, 28702800.0, 28706400.0, 28710000.0, 28713600.0, 28717200.0, 28720800.0, 28724400.0, 28728000.0, 28731600.0, 28735200.0, 28738800.0, 28742400.0, 28746000.0, 28749600.0, 28753200.0, 28756800.0, 28760400.0, 28764000.0, 28767600.0, 28771200.0, 28774800.0, 28778400.0, 28782000.0, 28785600.0, 28789200.0, 28792800.0, 28796400.0, 28800000.0, 28803600.0, 28807200.0, 28810800.0, 28814400.0, 28818000.0, 28821600.0, 28825200.0, 28828800.0, 28832400.0, 28836000.0, 28839600.0, 28843200.0, 28846800.0, 28850400.0, 28854000.0, 28857600.0, 28861200.0, 28864800.0, 28868400.0, 28872000.0, 28875600.0, 28879200.0, 28882800.0, 28886400.0, 28890000.0, 28893600.0, 28897200.0, 28900800.0, 28904400.0, 28908000.0, 28911600.0, 28915200.0, 28918800.0, 28922400.0, 28926000.0, 28929600.0, 28933200.0, 28936800.0, 28940400.0, 28944000.0, 28947600.0, 28951200.0, 28954800.0, 28958400.0, 28962000.0, 28965600.0, 28969200.0, 28972800.0, 28976400.0, 28980000.0, 28983600.0, 28987200.0, 28990800.0, 28994400.0, 28998000.0, 29001600.0, 29005200.0, 29008800.0, 29012400.0, 29016000.0, 29019600.0, 29023200.0, 29026800.0, 29030400.0, 29034000.0, 29037600.0, 29041200.0, 29044800.0, 29048400.0, 29052000.0, 29055600.0, 29059200.0, 29062800.0, 29066400.0, 29070000.0, 29073600.0, 29077200.0, 29080800.0, 29084400.0, 29088000.0, 29091600.0, 29095200.0, 29098800.0, 29102400.0, 29106000.0, 29109600.0, 29113200.0, 29116800.0, 29120400.0, 29124000.0, 29127600.0, 29131200.0, 29134800.0, 29138400.0, 29142000.0, 29145600.0, 29149200.0, 29152800.0, 29156400.0, 29160000.0, 29163600.0, 29167200.0, 29170800.0, 29174400.0, 29178000.0, 29181600.0, 29185200.0, 29188800.0, 29192400.0, 29196000.0, 29199600.0, 29203200.0, 29206800.0, 29210400.0, 29214000.0, 29217600.0, 29221200.0, 29224800.0, 29228400.0, 29232000.0, 29235600.0, 29239200.0, 29242800.0, 29246400.0, 29250000.0, 29253600.0, 29257200.0, 29260800.0, 29264400.0, 29268000.0, 29271600.0, 29275200.0, 29278800.0, 29282400.0, 29286000.0, 29289600.0, 29293200.0, 29296800.0, 29300400.0, 29304000.0, 29307600.0, 29311200.0, 29314800.0, 29318400.0, 29322000.0, 29325600.0, 29329200.0, 29332800.0, 29336400.0, 29340000.0, 29343600.0, 29347200.0, 29350800.0, 29354400.0, 29358000.0, 29361600.0, 29365200.0, 29368800.0, 29372400.0, 29376000.0, 29379600.0, 29383200.0, 29386800.0, 29390400.0, 29394000.0, 29397600.0, 29401200.0, 29404800.0, 29408400.0, 29412000.0, 29415600.0, 29419200.0, 29422800.0, 29426400.0, 29430000.0, 29433600.0, 29437200.0, 29440800.0, 29444400.0, 29448000.0, 29451600.0, 29455200.0, 29458800.0, 29462400.0, 29466000.0, 29469600.0, 29473200.0, 29476800.0, 29480400.0, 29484000.0, 29487600.0, 29491200.0, 29494800.0, 29498400.0, 29502000.0, 29505600.0, 29509200.0, 29512800.0, 29516400.0, 29520000.0, 29523600.0, 29527200.0, 29530800.0, 29534400.0, 29538000.0, 29541600.0, 29545200.0, 29548800.0, 29552400.0, 29556000.0, 29559600.0, 29563200.0, 29566800.0, 29570400.0, 29574000.0, 29577600.0, 29581200.0, 29584800.0, 29588400.0, 29592000.0, 29595600.0, 29599200.0, 29602800.0, 29606400.0, 29610000.0, 29613600.0, 29617200.0, 29620800.0, 29624400.0, 29628000.0, 29631600.0, 29635200.0, 29638800.0, 29642400.0, 29646000.0, 29649600.0, 29653200.0, 29656800.0, 29660400.0, 29664000.0, 29667600.0, 29671200.0, 29674800.0, 29678400.0, 29682000.0, 29685600.0, 29689200.0, 29692800.0, 29696400.0, 29700000.0, 29703600.0, 29707200.0, 29710800.0, 29714400.0, 29718000.0, 29721600.0, 29725200.0, 29728800.0, 29732400.0, 29736000.0, 29739600.0, 29743200.0, 29746800.0, 29750400.0, 29754000.0, 29757600.0, 29761200.0, 29764800.0, 29768400.0, 29772000.0, 29775600.0, 29779200.0, 29782800.0, 29786400.0, 29790000.0, 29793600.0, 29797200.0, 29800800.0, 29804400.0, 29808000.0, 29811600.0, 29815200.0, 29818800.0, 29822400.0, 29826000.0, 29829600.0, 29833200.0, 29836800.0, 29840400.0, 29844000.0, 29847600.0, 29851200.0, 29854800.0, 29858400.0, 29862000.0, 29865600.0, 29869200.0, 29872800.0, 29876400.0, 29880000.0, 29883600.0, 29887200.0, 29890800.0, 29894400.0, 29898000.0, 29901600.0, 29905200.0, 29908800.0, 29912400.0, 29916000.0, 29919600.0, 29923200.0, 29926800.0, 29930400.0, 29934000.0, 29937600.0, 29941200.0, 29944800.0, 29948400.0, 29952000.0, 29955600.0, 29959200.0, 29962800.0, 29966400.0, 29970000.0, 29973600.0, 29977200.0, 29980800.0, 29984400.0, 29988000.0, 29991600.0, 29995200.0, 29998800.0, 30002400.0, 30006000.0, 30009600.0, 30013200.0, 30016800.0, 30020400.0, 30024000.0, 30027600.0, 30031200.0, 30034800.0, 30038400.0, 30042000.0, 30045600.0, 30049200.0, 30052800.0, 30056400.0, 30060000.0, 30063600.0, 30067200.0, 30070800.0, 30074400.0, 30078000.0, 30081600.0, 30085200.0, 30088800.0, 30092400.0, 30096000.0, 30099600.0, 30103200.0, 30106800.0, 30110400.0, 30114000.0, 30117600.0, 30121200.0, 30124800.0, 30128400.0, 30132000.0, 30135600.0, 30139200.0, 30142800.0, 30146400.0, 30150000.0, 30153600.0, 30157200.0, 30160800.0, 30164400.0, 30168000.0, 30171600.0, 30175200.0, 30178800.0, 30182400.0, 30186000.0, 30189600.0, 30193200.0, 30196800.0, 30200400.0, 30204000.0, 30207600.0, 30211200.0, 30214800.0, 30218400.0, 30222000.0, 30225600.0, 30229200.0, 30232800.0, 30236400.0, 30240000.0, 30243600.0, 30247200.0, 30250800.0, 30254400.0, 30258000.0, 30261600.0, 30265200.0, 30268800.0, 30272400.0, 30276000.0, 30279600.0, 30283200.0, 30286800.0, 30290400.0, 30294000.0, 30297600.0, 30301200.0, 30304800.0, 30308400.0, 30312000.0, 30315600.0, 30319200.0, 30322800.0, 30326400.0, 30330000.0, 30333600.0, 30337200.0, 30340800.0, 30344400.0, 30348000.0, 30351600.0, 30355200.0, 30358800.0, 30362400.0, 30366000.0, 30369600.0, 30373200.0, 30376800.0, 30380400.0, 30384000.0, 30387600.0, 30391200.0, 30394800.0, 30398400.0, 30402000.0, 30405600.0, 30409200.0, 30412800.0, 30416400.0, 30420000.0, 30423600.0, 30427200.0, 30430800.0, 30434400.0, 30438000.0, 30441600.0, 30445200.0, 30448800.0, 30452400.0, 30456000.0, 30459600.0, 30463200.0, 30466800.0, 30470400.0, 30474000.0, 30477600.0, 30481200.0, 30484800.0, 30488400.0, 30492000.0, 30495600.0, 30499200.0, 30502800.0, 30506400.0, 30510000.0, 30513600.0, 30517200.0, 30520800.0, 30524400.0, 30528000.0, 30531600.0, 30535200.0, 30538800.0, 30542400.0, 30546000.0, 30549600.0, 30553200.0, 30556800.0, 30560400.0, 30564000.0, 30567600.0, 30571200.0, 30574800.0, 30578400.0, 30582000.0, 30585600.0, 30589200.0, 30592800.0, 30596400.0, 30600000.0, 30603600.0, 30607200.0, 30610800.0, 30614400.0, 30618000.0, 30621600.0, 30625200.0, 30628800.0, 30632400.0, 30636000.0, 30639600.0, 30643200.0, 30646800.0, 30650400.0, 30654000.0, 30657600.0, 30661200.0, 30664800.0, 30668400.0, 30672000.0, 30675600.0, 30679200.0, 30682800.0, 30686400.0, 30690000.0, 30693600.0, 30697200.0, 30700800.0, 30704400.0, 30708000.0, 30711600.0, 30715200.0, 30718800.0, 30722400.0, 30726000.0, 30729600.0, 30733200.0, 30736800.0, 30740400.0, 30744000.0, 30747600.0, 30751200.0, 30754800.0, 30758400.0, 30762000.0, 30765600.0, 30769200.0, 30772800.0, 30776400.0, 30780000.0, 30783600.0, 30787200.0, 30790800.0, 30794400.0, 30798000.0, 30801600.0, 30805200.0, 30808800.0, 30812400.0, 30816000.0, 30819600.0, 30823200.0, 30826800.0, 30830400.0, 30834000.0, 30837600.0, 30841200.0, 30844800.0, 30848400.0, 30852000.0, 30855600.0, 30859200.0, 30862800.0, 30866400.0, 30870000.0, 30873600.0, 30877200.0, 30880800.0, 30884400.0, 30888000.0, 30891600.0, 30895200.0, 30898800.0, 30902400.0, 30906000.0, 30909600.0, 30913200.0, 30916800.0, 30920400.0, 30924000.0, 30927600.0, 30931200.0, 30934800.0, 30938400.0, 30942000.0, 30945600.0, 30949200.0, 30952800.0, 30956400.0, 30960000.0, 30963600.0, 30967200.0, 30970800.0, 30974400.0, 30978000.0, 30981600.0, 30985200.0, 30988800.0, 30992400.0, 30996000.0, 30999600.0, 31003200.0, 31006800.0, 31010400.0, 31014000.0, 31017600.0, 31021200.0, 31024800.0, 31028400.0, 31032000.0, 31035600.0, 31039200.0, 31042800.0, 31046400.0, 31050000.0, 31053600.0, 31057200.0, 31060800.0, 31064400.0, 31068000.0, 31071600.0, 31075200.0, 31078800.0, 31082400.0, 31086000.0, 31089600.0, 31093200.0, 31096800.0, 31100400.0, 31104000.0, 31107600.0, 31111200.0, 31114800.0, 31118400.0, 31122000.0, 31125600.0, 31129200.0, 31132800.0, 31136400.0, 31140000.0, 31143600.0, 31147200.0, 31150800.0, 31154400.0, 31158000.0, 31161600.0, 31165200.0, 31168800.0, 31172400.0, 31176000.0, 31179600.0, 31183200.0, 31186800.0, 31190400.0, 31194000.0, 31197600.0, 31201200.0, 31204800.0, 31208400.0, 31212000.0, 31215600.0, 31219200.0, 31222800.0, 31226400.0, 31230000.0, 31233600.0, 31237200.0, 31240800.0, 31244400.0, 31248000.0, 31251600.0, 31255200.0, 31258800.0, 31262400.0, 31266000.0, 31269600.0, 31273200.0, 31276800.0, 31280400.0, 31284000.0, 31287600.0, 31291200.0, 31294800.0, 31298400.0, 31302000.0, 31305600.0, 31309200.0, 31312800.0, 31316400.0, 31320000.0, 31323600.0, 31327200.0, 31330800.0, 31334400.0, 31338000.0, 31341600.0, 31345200.0, 31348800.0, 31352400.0, 31356000.0, 31359600.0, 31363200.0, 31366800.0, 31370400.0, 31374000.0, 31377600.0, 31381200.0, 31384800.0, 31388400.0, 31392000.0, 31395600.0, 31399200.0, 31402800.0, 31406400.0, 31410000.0, 31413600.0, 31417200.0, 31420800.0, 31424400.0, 31428000.0, 31431600.0, 31435200.0, 31438800.0, 31442400.0, 31446000.0, 31449600.0, 31453200.0, 31456800.0, 31460400.0, 31464000.0, 31467600.0, 31471200.0, 31474800.0, 31478400.0, 31482000.0, 31485600.0, 31489200.0, 31492800.0, 31496400.0, 31500000.0, 31503600.0, 31507200.0, 31510800.0, 31514400.0, 31518000.0, 31521600.0, 31525200.0, 31528800.0, 31532400.0, 31536000.0;
     temp_year=
        7.9, 6.5, 5.2, 4.4, 4.4, 4.4, 4.1, 3.9, 3.1, 2.8, 3.5, 3.8, 4.2, 4.1, 4.2, 2.3, 3.3, 3.1, 2.9, 2.1, 1.7, 1.5, 1.3, 1.2, 0.7, 0.6, 1.2, 1.0, 0.8, 0.3, 0.2, 0.3, 1.0, 0.4, 2.0, 2.0, 2.2, 2.1, 2.2, 2.2, 2.3, 1.7, 1.9, 2.1, 2.0, 1.4, 1.2, 0.8, 0.6, 0.6, 0.6, 0.2, 0.3, -0.1, -0.1, 0.0, -0.2, -0.3, 0.1, 0.6, 1.4, 2.0, 2.1, 1.8, 0.4, -0.3, -1.2, -1.6, -1.2, -0.8, -1.3, -1.5, -2.8, -3.1, -3.6, -3.7, -4.2, -4.8, -5.2, -5.6, -6.1, -6.1, -4.5, -3.2, -2.0, -1.1, -0.4, -0.5, -0.9, -1.5, -2.9, -3.4, -4.1, -4.7, -5.4, -5.9, -5.9, -6.1, -6.2, -6.4, -6.2, -6.7, -6.5, -7.0, -6.9, -7.0, -6.2, -4.3, -2.9, -2.9, -1.8, -2.9, -2.9, -3.8, -4.9, -6.0, -6.9, -6.8, -6.5, -7.1, -7.2, -6.8, -7.3, -7.0, -7.6, -7.5, -7.3, -8.3, -9.1, -9.3, -7.4, -4.9, -4.4, -3.3, -3.3, -3.4, -3.6, -4.2, -5.2, -6.4, -7.4, -8.0, -7.3, -5.7, -5.1, -4.9, -4.9, -4.5, -4.3, -4.2, -4.0, -3.9, -3.6, -3.5, -3.3, -3.1, -2.6, -2.2, -2.0, -1.9, -2.1, -2.3, -2.3, -2.5, -3.0, -3.3, -3.6, -3.8, -3.9, -3.9, -3.9, -3.9, -4.2, -4.5, -4.7, -4.9, -5.0, -5.1, -5.1, -4.6, -3.4, -2.6, -2.4, -1.9, -1.9, -2.2, -2.6, -2.8, -2.8, -3.2, -3.1, -2.5, -2.2, -2.4, -3.0, -2.8, -2.8, -2.6, -2.5, -2.3, -2.0, -1.7, -1.4, -0.9, -0.3, 0.1, 0.4, 0.8, 0.9, 1.1, 1.1, 1.3, 1.1, 1.1, 1.3, 1.1, 1.2, 1.4, 2.1, 2.7, 3.4, 3.5, 3.7, 3.8, 4.4, 5.4, 5.6, 6.0, 6.9, 7.1, 6.5, 6.6, 6.0, 5.1, 4.7, 4.4, 4.4, 4.5, 3.4, 2.9, 2.1, 1.7, 2.0, 2.8, 3.1, 4.8, 3.2, 3.2, 3.3, 2.9, 2.7, 3.8, 2.9, 3.4, 3.6, 3.7, 3.9, 3.7, 3.1, 3.1, 3.0, 2.7, 2.8, 2.6, 2.7, 2.7, 2.1, 2.5, 2.4, 2.2, 2.1, 2.3, 2.1, 1.5, 1.7, 0.9, 0.5, 1.2, 1.9, 2.9, 2.8, 2.2, 1.8, 1.5, 0.9, 0.7, 0.5, 0.7, 0.4, 0.2, -0.3, -0.5, -1.7, -3.0, -3.2, -4.1, -3.7, -2.8, -2.2, 0.0, 1.7, 2.0, 2.5, 1.3, 1.0, -0.4, -2.2, -3.0, -2.7, -2.9, -2.2, -1.4, -2.4, -2.7, -2.7, -2.7, -2.8, -2.7, -2.4, -2.1, -2.2, -2.1, -1.9, -1.6, -1.4, -0.8, -0.2, -0.2, 0.1, -0.3, -0.3, -0.2, -0.2, -0.2, -0.6, -0.6, -0.6, -0.4, -0.4, -0.2, -0.1, -0.1, -0.1, 0.1, 0.2, 0.3, 0.5, 0.8, 1.2, 1.6, 1.7, 2.1, 2.1, 1.9, 1.8, 1.9, 1.8, 1.7, 1.6, 1.7, 1.4, 1.8, 2.1, 2.0, 1.7, 1.4, 1.4, 1.4, 1.6, 0.8, 1.8, 3.9, 4.0, 5.7, 5.9, 3.8, 3.6, 1.3, -0.4, -0.4, -0.8, -1.1, -1.1, -1.4, -1.5, -2.0, -2.5, -2.9, -3.4, -3.4, -3.8, -4.3, -4.5, -4.9, -2.5, -0.8, 1.5, 3.6, 5.1, 4.0, 4.4, 2.6, 0.1, -0.7, -1.5, -1.9, -2.6, -3.0, -3.8, -3.7, -3.7, -3.8, -3.8, -3.5, -3.4, -3.0, -2.2, -1.8, -1.0, -0.4, 0.0, 0.2, 0.4, 0.3, 0.5, 0.6, 0.7, 0.8, 0.6, 0.5, 0.8, 0.7, 1.0, 1.2, 1.1, 1.3, 1.6, 1.6, 1.6, 1.8, 1.8, 2.0, 1.5, 2.7, 5.0, 6.8, 6.5, 6.5, 6.7, 5.0, 3.3, 2.9, 3.3, 3.8, 3.1, 2.5, 3.1, 3.2, 3.2, 3.3, 3.9, 3.5, 2.9, 2.4, 1.2, 1.8, 3.2, 3.6, 4.0, 3.9, 5.0, 5.4, 5.5, 5.1, 4.6, 4.8, 4.2, 5.0, 4.3, 4.3, 4.5, 4.5, 4.2, 4.0, 3.4, 3.2, 3.1, 3.0, 2.9, 3.0, 3.6, 5.3, 5.9, 6.2, 7.1, 7.3, 6.8, 6.0, 4.8, 5.7, 5.0, 5.5, 5.9, 6.3, 7.0, 7.0, 6.3, 6.1, 6.1, 6.2, 6.5, 6.9, 7.9, 7.6, 8.2, 8.0, 8.7, 8.7, 8.5, 8.6, 8.9, 9.4, 9.9, 10.9, 10.6, 10.6, 10.9, 12.3, 12.6, 12.9, 12.7, 11.8, 11.8, 11.2, 10.8, 10.8, 8.9, 8.7, 8.0, 7.8, 8.0, 7.9, 8.1, 8.1, 7.9, 7.6, 6.5, 6.1, 5.6, 5.7, 5.9, 6.5, 6.8, 6.7, 6.5, 6.0, 5.8, 4.3, 4.0, 4.7, 5.1, 5.4, 5.7, 6.1, 7.0, 6.1, 5.6, 6.3, 6.6, 6.6, 6.4, 5.9, 5.8, 4.8, 5.2, 4.9, 5.0, 4.5, 4.4, 4.2, 4.1, 4.3, 3.4, 1.7, 2.7, 3.3, 4.0, 5.0, 6.3, 9.6, 10.5, 10.8, 11.1, 12.5, 12.4, 11.3, 11.9, 11.8, 11.8, 11.6, 11.0, 11.5, 11.8, 11.9, 12.2, 12.1, 11.7, 12.1, 10.7, 11.0, 12.1, 13.4, 12.9, 13.4, 13.1, 13.2, 11.9, 11.0, 11.5, 8.0, 7.5, 7.1, 6.1, 3.5, 3.7, 3.7, 3.4, 3.1, 3.0, 2.6, 1.6, 1.3, 1.5, 1.7, 2.9, 3.1, 3.5, 4.1, 4.9, 5.0, 4.8, 3.7, 2.4, 2.4, 2.1, 2.5, 2.6, 3.0, 3.5, 3.8, 4.1, 4.5, 4.4, 4.4, 4.7, 5.4, 5.8, 6.0, 6.7, 8.8, 9.4, 10.3, 10.2, 10.4, 8.9, 9.1, 6.5, 6.3, 6.8, 6.4, 6.3, 6.6, 6.9, 6.7, 7.4, 8.0, 7.3, 6.6, 6.5, 6.4, 7.0, 7.7, 8.3, 9.9, 9.6, 9.2, 8.3, 8.4, 8.5, 8.8, 8.5, 8.4, 9.6, 10.0, 9.5, 9.1, 9.3, 8.0, 8.1, 8.0, 7.8, 7.8, 7.7, 7.5, 7.6, 7.8, 8.4, 7.5, 7.4, 7.2, 5.9, 5.5, 4.9, 4.5, 4.0, 3.2, 1.8, 0.8, -0.2, 0.5, 2.0, 4.1, 5.9, 7.2, 7.2, 7.2, 6.9, 9.2, 9.1, 9.2, 9.3, 9.8, 12.0, 14.0, 13.9, 13.8, 13.7, 12.0, 9.4, 9.2, 6.9, 6.6, 4.7, 5.8, 5.8, 7.6, 8.2, 7.4, 7.6, 5.9, 6.1, 6.6, 7.7, 8.5, 9.4, 10.2, 10.3, 10.8, 11.1, 11.9, 11.7, 11.4, 11.2, 10.9, 11.1, 10.5, 9.8, 9.4, 8.2, 8.6, 9.2, 7.5, 7.9, 8.5, 7.1, 7.6, 7.0, 8.1, 11.1, 12.3, 13.3, 15.2, 16.0, 16.8, 16.4, 15.2, 10.8, 8.6, 7.6, 7.6, 5.6, 4.3, 3.9, 4.7, 3.7, 2.8, 2.2, 1.3, 1.2, 1.5, 2.3, 3.5, 7.9, 11.1, 13.0, 13.9, 14.4, 14.6, 15.2, 13.6, 9.8, 7.2, 6.9, 5.9, 4.0, 4.2, 3.8, 4.4, 6.3, 10.4, 11.1, 11.5, 10.5, 9.3, 8.3, 7.3, 9.1, 10.8, 12.3, 11.9, 12.6, 12.5, 12.2, 10.2, 7.0, 6.0, 7.7, 8.4, 8.9, 8.4, 9.6, 9.5, 10.1, 9.5, 9.6, 10.8, 11.7, 11.6, 11.8, 12.4, 13.5, 13.5, 13.6, 15.3, 15.3, 15.4, 13.4, 13.7, 13.0, 12.0, 10.9, 10.3, 10.0, 9.7, 8.8, 8.8, 8.2, 8.1, 8.4, 8.6, 7.6, 8.6, 8.0, 8.4, 8.8, 9.2, 9.6, 10.1, 10.3, 10.3, 10.0, 9.6, 9.1, 8.9, 7.5, 7.6, 7.8, 6.8, 6.0, 5.4, 4.4, 4.4, 2.5, 1.7, 1.5, 1.4, 2.5, 3.6, 4.6, 5.6, 6.5, 8.7, 10.4, 9.5, 9.1, 7.9, 7.4, 7.0, 6.7, 6.2, 5.8, 5.4, 5.7, 6.5, 5.7, 4.9, 4.7, 4.7, 4.9, 5.0, 5.4, 5.6, 6.5, 6.9, 6.9, 6.9, 7.0, 7.1, 7.3, 7.5, 7.3, 7.0, 7.1, 7.4, 7.3, 7.6, 7.7, 8.1, 8.2, 8.5, 8.6, 8.7, 9.0, 9.3, 9.5, 9.8, 10.3, 11.2, 11.4, 12.3, 12.4, 12.0, 12.1, 12.0, 11.6, 10.2, 10.2, 9.6, 9.1, 7.0, 4.4, 1.2, -0.9, -2.2, -1.5, -1.0, 0.5, 0.7, 0.8, 1.0, 1.5, 1.9, 2.3, 3.2, 3.5, 3.8, 3.7, 3.3, 2.9, 2.6, 2.4, 0.9, 2.2, 2.1, 1.9, 1.9, 1.7, 1.6, 1.4, 1.3, 1.3, 1.3, 1.2, 1.1, 1.4, 1.6, 1.9, 2.0, 2.1, 2.3, 2.8, 2.8, 2.0, 0.9, -0.3, -0.7, -1.0, -1.6, -2.2, -2.7, -3.5, -4.2, -3.9, -3.2, -2.2, -1.9, -1.8, -1.3, -0.9, -0.5, 0.2, 0.8, 0.9, 1.1, 1.0, 0.9, 0.6, 0.6, 0.4, 0.4, 0.4, 0.4, 0.4, 0.0, -0.1, -0.2, -0.4, -0.6, -0.7, -0.8, -0.7, -0.7, -0.7, -0.5, -0.5, -0.3, -0.2, 0.1, 0.4, 0.4, 0.2, 0.2, 0.1, 0.2, 0.2, 0.2, 0.1, -0.1, -0.1, -0.2, -0.9, -1.0, -1.2, -1.2, -1.3, -1.3, -1.3, -1.0, -0.9, -0.2, 0.1, 0.7, 1.5, 0.6, -0.1, -0.2, -0.4, -0.1, 0.0, -0.2, -0.3, -0.4, -0.6, -0.7, -1.3, -1.3, -1.1, -1.1, -0.9, -1.1, -1.0, -0.9, -0.7, -0.7, -0.5, -0.1, 0.0, -0.2, -0.3, -0.3, -0.5, -0.5, -0.6, -0.7, -0.8, -0.8, -0.9, -1.0, -1.1, -1.0, -1.6, -1.7, -1.5, -1.6, -1.3, -1.1, -0.3, 0.1, 0.5, 0.8, 0.9, 1.2, 1.0, 1.0, 0.7, 0.7, 0.8, 0.8, 0.8, 0.9, 0.9, 0.8, 0.8, 0.5, 0.5, 0.5, 0.7, 0.7, 0.7, 0.9, 1.4, 1.5, 2.0, 2.4, 2.8, 2.8, 3.1, 3.1, 3.1, 3.0, 3.1, 2.8, 2.7, 2.9, 2.8, 2.6, 2.5, 2.4, 2.4, 2.2, 2.3, 2.7, 3.8, 4.4, 5.3, 5.6, 6.4, 6.6, 6.5, 6.5, 6.1, 5.6, 3.7, 3.1, 3.8, 4.3, 4.0, 4.0, 3.9, 3.7, 4.6, 4.4, 4.2, 4.2, 5.0, 5.1, 6.0, 6.6, 6.7, 6.4, 7.3, 7.0, 6.0, 6.3, 6.4, 5.0, 4.9, 4.0, 4.0, 4.3, 4.2, 4.8, 4.8, 4.6, 3.9, 3.8, 4.0, 3.7, 4.3, 3.9, 3.9, 4.2, 4.9, 5.0, 5.8, 6.7, 6.6, 6.3, 5.7, 5.4, 5.4, 5.1, 5.8, 6.0, 6.0, 5.7, 4.7, 4.9, 4.8, 2.3, 2.3, 2.8, 2.8, 1.9, 3.4, 3.6, 3.6, 4.8, 5.4, 6.2, 5.8, 4.9, 4.2, 3.5, 1.3, 1.3, 1.8, 1.8, 1.4, 0.8, 0.4, 0.1, -0.3, -0.7, -1.1, -1.8, -2.5, -0.5, 0.7, 1.6, 1.8, 2.6, 3.1, 3.7, 3.2, 2.2, 1.1, -0.3, -2.5, -3.7, -4.2, -5.8, -5.1, -5.8, -6.0, -6.1, -5.4, -7.0, -6.8, -5.3, -3.8, -2.7, -2.0, -1.2, -1.4, -0.4, -0.2, -0.8, -1.1, -1.4, -1.7, -2.8, -3.7, -3.6, -3.9, -5.4, -6.6, -6.6, -6.7, -6.8, -7.9, -8.2, -8.6, -8.6, -8.6, -6.1, -3.9, -1.2, -0.5, 0.4, 1.4, 2.5, 2.2, 1.3, 0.6, -0.6, -3.9, -3.5, -3.4, -3.6, -5.5, -5.2, -5.5, -5.9, -7.2, -8.5, -8.9, -9.0, -8.8, -6.2, -4.3, -1.8, -0.2, 0.5, 1.9, 2.2, 3.4, 1.7, 0.6, -0.3, -0.7, -1.3, -1.8, -2.5, -3.3, -3.9, -4.4, -4.7, -4.8, -4.6, -4.8, -4.9, -2.0, 1.1, 2.5, 3.8, 4.6, 7.4, 9.9, 11.8, 12.8, 12.4, 10.1, 7.5, 3.8, 3.7, 3.9, 3.5, 1.0, 2.3, -0.5, -1.9, -2.6, -3.2, -3.3, -4.2, -3.6, -0.2, 4.0, 5.6, 7.8, 8.3, 9.0, 10.1, 12.1, 12.0, 10.0, 7.2, 4.2, 4.2, 2.6, 1.7, -0.3, 0.0, 1.3, 1.4, 1.7, 3.7, 4.1, 4.1, 4.2, 6.1, 8.5, 10.5, 12.3, 13.8, 13.7, 14.0, 14.2, 13.7, 10.4, 8.7, 8.4, 7.5, 6.5, 6.1, 5.5, 6.8, 6.2, 7.0, 7.4, 6.1, 6.1, 6.0, 6.0, 6.6, 7.7, 7.8, 8.7, 9.1, 9.9, 10.8, 11.5, 11.2, 9.8, 9.5, 9.1, 8.9, 8.3, 8.5, 7.6, 7.2, 7.9, 7.8, 7.9, 7.6, 7.5, 7.5, 7.4, 7.7, 10.2, 11.6, 11.6, 11.1, 10.5, 8.5, 8.9, 9.1, 8.4, 7.6, 6.8, 6.4, 6.1, 6.1, 6.0, 6.0, 6.0, 5.6, 5.3, 5.3, 5.5, 5.2, 5.5, 5.5, 5.6, 5.9, 6.5, 6.9, 7.1, 7.5, 7.1, 6.9, 6.5, 6.3, 6.3, 6.1, 5.8, 5.3, 4.9, 4.5, 2.8, 1.3, 2.6, 3.3, 3.7, 3.9, 4.1, 5.6, 7.8, 8.9, 9.0, 10.2, 10.3, 11.1, 11.4, 10.3, 9.3, 7.8, 6.8, 6.1, 5.9, 5.9, 6.1, 6.1, 6.1, 6.6, 6.3, 6.5, 6.3, 6.9, 6.7, 7.8, 8.0, 9.6, 9.7, 10.8, 12.3, 13.2, 14.1, 13.9, 13.0, 11.4, 10.8, 10.1, 10.7, 9.7, 8.6, 6.8, 7.3, 7.7, 7.3, 5.9, 6.7, 5.9, 5.1, 7.1, 8.5, 9.7, 9.7, 9.6, 8.4, 7.5, 8.5, 7.2, 6.5, 6.5, 6.4, 6.2, 6.2, 6.0, 5.5, 5.2, 4.8, 3.0, 1.3, 1.0, 0.3, 0.3, 0.7, 3.3, 6.0, 8.1, 8.8, 9.4, 10.2, 10.4, 11.0, 9.9, 8.2, 6.7, 6.4, 6.2, 6.1, 5.5, 4.6, 3.3, 2.2, 1.3, 1.0, 0.7, 0.6, -0.4, 0.2, 2.8, 4.7, 4.7, 6.2, 6.0, 6.5, 7.4, 7.3, 6.5, 5.1, 3.7, 2.8, 2.3, 1.2, 1.1, 0.3, 0.1, -0.7, -1.2, -0.7, -0.9, -1.4, -1.8, -2.4, 0.8, 3.0, 4.6, 6.2, 6.8, 7.7, 8.0, 8.0, 7.0, 5.4, 3.0, 1.4, -0.8, -1.5, -2.5, -2.9, -2.8, -3.0, -3.1, -3.8, -4.1, -2.9, -1.8, -1.0, 2.6, 5.0, 6.7, 9.0, 11.1, 14.0, 13.7, 13.2, 12.0, 10.3, 9.2, 8.2, 7.0, 7.0, 6.4, 5.7, 5.7, 5.4, 5.3, 5.4, 5.3, 5.3, 5.2, 5.5, 6.7, 7.8, 8.0, 8.9, 10.4, 11.6, 12.5, 12.9, 12.8, 11.8, 10.1, 8.1, 6.0, 5.3, 3.6, 2.7, 1.1, 0.5, -0.4, -0.2, -0.1, -1.6, -1.9, -1.7, 2.9, 8.5, 10.9, 12.4, 14.0, 15.2, 16.6, 16.8, 16.4, 13.9, 10.2, 8.2, 6.5, 5.6, 2.9, 2.2, 2.5, 2.3, 0.3, -0.1, -1.0, -1.3, -1.2, -0.7, 4.8, 8.2, 11.8, 13.0, 13.9, 16.1, 17.0, 15.8, 16.3, 14.1, 11.4, 8.5, 6.3, 3.9, 2.6, 2.1, 0.8, 0.5, 0.2, -0.1, -0.4, 1.7, 1.7, 1.9, 7.3, 10.0, 12.3, 15.1, 15.7, 16.5, 17.4, 17.3, 17.1, 14.3, 12.0, 9.4, 7.1, 5.7, 3.6, 2.8, 2.9, 2.5, 2.1, 0.2, 0.0, -0.9, -1.1, 1.2, 6.0, 9.8, 11.5, 13.8, 16.4, 18.0, 19.0, 18.8, 17.5, 15.2, 11.8, 8.6, 6.2, 5.5, 5.0, 3.9, 3.8, 3.0, 2.2, 1.8, 3.1, 3.4, 5.4, 7.0, 7.5, 10.7, 15.1, 17.8, 18.9, 18.5, 19.9, 18.6, 17.5, 17.2, 16.5, 15.5, 15.2, 15.1, 15.6, 14.7, 13.8, 13.3, 13.0, 12.8, 12.4, 11.5, 10.4, 10.0, 10.0, 10.1, 9.8, 10.3, 10.7, 11.7, 12.1, 12.1, 13.1, 13.6, 13.5, 13.2, 11.6, 10.7, 8.8, 8.0, 7.2, 6.2, 5.3, 6.5, 8.3, 8.3, 8.2, 9.4, 11.2, 11.3, 11.4, 11.9, 12.8, 14.2, 15.0, 15.5, 15.8, 14.6, 13.5, 11.5, 12.8, 12.4, 12.0, 11.1, 10.3, 9.2, 8.1, 9.9, 9.9, 9.2, 8.6, 8.5, 9.9, 11.1, 11.5, 12.6, 14.1, 14.3, 14.8, 15.0, 15.0, 13.9, 13.0, 9.2, 5.8, 5.6, 4.5, 5.0, 4.8, 5.0, 4.5, 2.5, 0.6, 0.6, 0.7, 2.2, 4.2, 7.3, 9.9, 12.9, 13.9, 16.4, 17.4, 16.8, 17.1, 15.8, 14.2, 9.5, 7.0, 6.0, 4.6, 3.0, 3.1, 2.7, 2.3, 2.5, 2.1, 2.8, 2.6, 3.2, 8.3, 12.7, 14.7, 15.2, 14.8, 14.3, 14.2, 14.0, 13.7, 13.0, 12.1, 11.4, 1.1, 10.8, 10.9, 10.9, 9.7, 9.4, 9.0, 9.8, 10.1, 10.1, 10.2, 10.2, 11.0, 12.3, 13.8, 13.7, 13.5, 14.9, 14.1, 14.5, 13.6, 13.0, 13.0, 12.2, 11.8, 12.0, 11.7, 11.5, 11.4, 11.2, 11.0, 11.1, 10.8, 10.3, 9.7, 9.4, 9.5, 10.5, 12.1, 12.1, 12.3, 13.4, 13.0, 12.4, 11.8, 11.3, 10.5, 9.8, 9.7, 9.3, 8.8, 8.1, 7.4, 5.7, 5.2, 5.1, 4.5, 3.9, 4.2, 4.6, 5.7, 7.4, 8.7, 10.5, 10.6, 11.5, 10.4, 10.2, 9.8, 9.3, 8.6, 5.9, 4.7, 4.1, 3.2, 2.0, 1.0, 0.2, 0.0, -1.0, -1.5, -1.3, -0.3, 1.4, 4.8, 6.0, 6.7, 7.4, 8.3, 8.2, 6.7, 9.1, 8.8, 8.2, 7.1, 5.9, 4.7, 3.6, 2.6, 2.8, 2.9, 2.8, 2.7, 2.4, 2.4, 1.6, 1.0, 1.4, 3.7, 5.0, 6.6, 6.4, 8.2, 8.1, 8.8, 9.2, 7.6, 6.9, 5.0, 4.2, 2.5, 1.6, 0.8, 0.6, -1.0, -1.2, -2.2, -1.6, -1.2, -1.8, -2.2, -1.4, 1.3, 2.9, 4.6, 5.8, 6.0, 6.0, 5.6, 5.1, 5.0, 4.4, 3.5, 2.7, 1.5, 0.8, -0.1, -0.2, -0.5, -1.0, -1.2, -2.0, -3.0, -3.2, -2.8, -1.6, 1.2, 2.9, 5.0, 5.5, 6.4, 5.6, 6.2, 7.0, 6.4, 4.9, 3.8, 2.3, 1.3, -0.4, -2.0, -1.0, -1.9, -2.6, -2.8, -5.1, -6.2, -6.6, -5.3, -1.8, 1.1, 4.3, 5.4, 6.3, 7.7, 7.7, 7.8, 8.3, 7.8, 6.8, 5.0, 2.7, 0.9, -0.5, -1.3, -1.7, -1.7, -1.5, -1.4, -1.7, -1.9, -2.7, -1.6, 1.7, 4.6, 7.8, 10.0, 13.1, 13.2, 14.2, 15.8, 15.2, 14.8, 13.7, 11.7, 9.2, 7.1, 4.2, 6.7, 6.2, 5.1, 7.1, 6.3, 6.3, 6.2, 4.7, 6.4, 7.6, 9.3, 12.6, 13.9, 15.5, 16.9, 17.0, 17.8, 18.3, 18.0, 16.7, 14.8, 13.1, 11.6, 11.0, 10.4, 9.9, 8.5, 6.7, 6.0, 5.0, 6.6, 6.2, 6.3, 7.4, 8.5, 10.0, 12.0, 13.0, 14.9, 17.1, 18.1, 17.4, 17.8, 17.6, 15.7, 12.2, 10.2, 8.0, 5.7, 5.3, 5.0, 4.6, 3.0, 3.1, 4.4, 5.3, 5.2, 5.4, 9.6, 12.4, 15.0, 16.9, 18.8, 19.8, 21.5, 20.6, 20.3, 18.8, 17.0, 15.4, 14.8, 14.7, 14.9, 14.4, 11.6, 11.0, 8.4, 7.4, 5.9, 5.0, 6.7, 9.4, 11.7, 13.7, 15.2, 16.6, 18.0, 18.9, 19.6, 20.7, 19.7, 19.5, 18.1, 16.3, 16.1, 14.6, 12.9, 11.4, 12.0, 13.2, 13.3, 11.9, 12.7, 12.1, 11.8, 12.0, 12.6, 12.9, 14.1, 15.1, 16.6, 16.5, 16.8, 15.9, 15.7, 15.1, 14.6, 13.5, 10.5, 9.3, 7.0, 6.9, 6.5, 6.1, 7.9, 6.9, 7.3, 9.0, 9.3, 10.5, 11.4, 11.9, 12.5, 11.3, 11.7, 12.9, 14.4, 15.8, 15.7, 15.0, 14.0, 13.1, 10.1, 7.5, 7.5, 7.7, 8.2, 8.5, 8.5, 8.3, 8.2, 8.6, 7.9, 9.4, 10.0, 6.9, 9.3, 11.1, 10.9, 12.3, 12.8, 11.5, 9.8, 10.9, 9.5, 9.4, 9.5, 7.3, 7.1, 7.6, 7.6, 7.7, 7.3, 7.3, 7.0, 5.0, 4.9, 5.1, 5.7, 6.7, 7.5, 8.7, 8.6, 10.6, 10.5, 11.4, 11.0, 9.4, 7.1, 6.1, 6.1, 6.0, 4.5, 4.6, 3.8, 3.8, 4.3, 3.7, 4.1, 4.0, 5.4, 5.6, 6.4, 8.7, 8.7, 8.8, 7.6, 10.0, 9.5, 10.5, 8.0, 7.6, 7.9, 6.7, 6.4, 5.9, 5.7, 5.3, 4.9, 4.4, 4.0, 3.4, 2.9, 1.7, 1.1, 2.0, 5.5, 5.7, 6.2, 7.3, 7.7, 8.1, 8.6, 8.5, 8.7, 9.1, 8.1, 6.6, 5.4, 4.5, 4.8, 4.9, 4.6, 5.6, 5.7, 4.8, 4.8, 4.6, 4.8, 4.8, 5.2, 5.4, 6.1, 6.6, 7.0, 7.0, 7.3, 7.4, 7.7, 7.9, 7.7, 7.5, 7.5, 7.4, 7.3, 7.1, 6.9, 6.9, 6.8, 6.7, 6.7, 6.5, 6.6, 7.2, 8.0, 9.7, 10.4, 11.6, 12.3, 12.3, 13.8, 14.6, 14.9, 13.6, 12.4, 10.6, 9.0, 7.7, 6.8, 5.9, 5.1, 4.7, 3.2, 1.8, 1.4, 1.0, 1.8, 4.4, 6.1, 6.9, 8.4, 10.9, 13.7, 12.9, 14.9, 12.7, 14.2, 10.6, 10.2, 9.7, 9.4, 8.6, 9.2, 8.5, 8.1, 7.4, 6.9, 6.9, 7.1, 7.3, 7.6, 7.7, 8.6, 8.7, 9.3, 9.9, 11.1, 11.4, 11.6, 12.5, 11.0, 10.8, 10.3, 9.5, 8.8, 7.4, 5.9, 4.7, 4.1, 3.2, 2.5, 1.8, 1.3, 1.3, 1.0, 5.5, 7.2, 8.5, 9.7, 11.6, 11.9, 12.7, 13.2, 13.5, 13.7, 13.7, 13.3, 12.8, 12.1, 10.3, 9.0, 7.7, 8.0, 6.5, 5.0, 2.8, 2.5, 1.7, 3.2, 5.9, 7.6, 9.6, 11.8, 13.4, 14.0, 14.6, 14.5, 14.6, 14.8, 14.3, 13.5, 12.5, 12.1, 9.8, 8.9, 8.4, 8.1, 8.2, 7.5, 7.1, 7.0, 6.6, 6.3, 7.0, 8.2, 9.6, 10.7, 8.6, 7.3, 10.3, 10.3, 11.1, 10.1, 10.1, 8.5, 8.0, 8.4, 8.5, 7.9, 7.7, 7.4, 7.3, 7.1, 7.0, 6.9, 6.8, 7.2, 7.6, 7.8, 8.6, 8.4, 9.1, 9.5, 9.4, 10.2, 10.5, 10.2, 9.7, 9.1, 8.8, 9.0, 9.3, 9.6, 9.1, 8.8, 8.4, 8.1, 8.4, 8.1, 8.0, 8.0, 8.5, 9.2, 9.5, 10.4, 10.8, 11.1, 11.2, 11.5, 11.3, 11.1, 11.5, 11.3, 10.6, 10.6, 10.4, 9.7, 9.0, 8.7, 8.4, 8.3, 8.4, 8.3, 7.9, 7.7, 7.3, 7.3, 7.7, 8.7, 9.5, 9.3, 9.8, 10.1, 10.3, 9.8, 8.7, 7.7, 7.2, 7.2, 6.9, 5.7, 4.9, 5.1, 5.2, 5.0, 4.9, 4.9, 4.6, 4.5, 4.6, 7.5, 7.6, 7.8, 7.9, 8.3, 9.2, 10.5, 10.6, 10.9, 10.1, 9.2, 7.7, 5.3, 5.0, 4.4, 4.0, 2.7, 2.7, 2.2, 2.1, 2.3, 3.6, 4.6, 6.1, 8.4, 9.9, 11.7, 12.7, 14.3, 13.7, 14.4, 14.7, 15.9, 16.1, 15.3, 14.6, 12.8, 13.5, 13.2, 12.7, 11.3, 10.4, 9.9, 8.8, 7.9, 7.6, 8.2, 8.1, 9.0, 10.5, 11.6, 12.9, 15.1, 15.8, 16.5, 17.0, 17.0, 15.7, 14.1, 13.3, 12.8, 11.5, 10.4, 9.2, 8.3, 9.0, 8.4, 8.0, 7.1, 6.5, 7.5, 10.2, 13.4, 15.6, 18.0, 19.7, 20.4, 21.7, 22.5, 22.8, 23.3, 22.9, 22.2, 20.6, 19.1, 18.3, 16.9, 16.3, 13.1, 13.3, 12.7, 12.1, 10.6, 10.4, 11.5, 14.2, 16.1, 17.5, 19.9, 21.4, 23.5, 25.5, 25.7, 25.5, 25.7, 25.2, 23.7, 22.2, 21.0, 20.1, 17.9, 15.6, 13.0, 11.1, 10.0, 10.4, 10.5, 11.1, 11.4, 11.0, 11.2, 11.5, 12.8, 14.8, 16.3, 19.1, 20.2, 18.7, 18.0, 17.4, 16.7, 16.1, 14.6, 14.4, 13.9, 13.3, 12.0, 11.5, 11.0, 10.9, 11.8, 12.1, 12.5, 12.5, 12.7, 13.9, 15.7, 17.0, 16.7, 17.4, 16.4, 16.2, 16.6, 16.0, 15.8, 15.0, 14.7, 14.0, 13.2, 12.9, 12.9, 13.3, 12.8, 13.0, 13.0, 12.2, 12.2, 12.7, 14.2, 16.2, 18.3, 18.8, 19.7, 20.3, 20.5, 20.2, 13.3, 12.8, 12.5, 11.3, 11.0, 10.6, 10.5, 10.3, 10.2, 10.0, 9.7, 9.3, 9.0, 9.1, 9.4, 9.8, 10.2, 10.7, 11.5, 11.7, 11.6, 12.2, 12.8, 12.4, 13.2, 12.9, 12.6, 11.8, 10.6, 9.3, 8.3, 7.4, 6.7, 6.8, 6.5, 5.9, 5.2, 4.6, 5.5, 8.0, 10.8, 12.5, 14.0, 13.8, 13.4, 13.1, 13.4, 13.4, 13.4, 13.2, 13.2, 12.8, 12.3, 12.1, 11.9, 11.8, 11.6, 11.1, 10.2, 8.4, 6.6, 6.8, 9.0, 12.9, 15.5, 16.9, 18.2, 20.4, 20.9, 21.2, 21.8, 22.1, 22.2, 20.5, 19.7, 18.1, 16.7, 15.8, 15.0, 14.1, 12.7, 12.2, 11.8, 11.3, 10.8, 11.1, 12.0, 13.4, 16.0, 18.4, 18.4, 19.0, 20.1, 21.2, 21.9, 21.7, 15.7, 11.9, 12.2, 12.3, 12.0, 12.0, 12.3, 12.5, 12.3, 11.6, 11.4, 11.5, 11.5, 11.6, 11.6, 12.2, 12.6, 13.6, 13.9, 13.6, 13.7, 13.9, 14.2, 14.5, 13.9, 13.8, 12.8, 12.5, 12.5, 12.3, 11.5, 11.2, 11.4, 11.2, 11.2, 11.2, 11.4, 11.4, 11.0, 10.9, 11.1, 11.1, 11.1, 12.0, 13.0, 13.1, 13.3, 13.8, 13.7, 13.1, 12.7, 12.1, 11.7, 11.3, 11.1, 10.9, 10.9, 10.8, 10.7, 10.5, 10.5, 10.3, 8.5, 9.3, 10.6, 11.0, 11.8, 11.3, 11.5, 13.0, 12.7, 12.5, 12.9, 12.9, 12.6, 10.9, 10.0, 9.1, 8.7, 8.5, 8.4, 8.2, 8.0, 7.5, 7.2, 6.4, 6.4, 6.9, 7.2, 7.4, 8.9, 8.7, 8.7, 9.1, 9.9, 9.5, 9.9, 9.7, 9.1, 7.9, 5.3, 4.3, 3.7, 3.2, 2.5, 2.6, 3.0, 2.4, 1.3, 1.9, 5.6, 9.2, 10.7, 11.0, 12.2, 12.8, 13.2, 13.2, 12.4, 11.1, 10.4, 10.7, 10.4, 10.3, 9.6, 8.1, 8.0, 7.5, 6.2, 5.6, 4.5, 4.6, 4.2, 4.4, 5.8, 7.7, 10.9, 13.2, 15.4, 18.3, 18.7, 19.6, 20.9, 20.9, 20.7, 20.6, 19.7, 17.6, 15.7, 16.4, 15.5, 14.5, 14.2, 13.9, 13.4, 13.6, 13.3, 13.6, 14.7, 15.0, 16.9, 18.2, 20.0, 21.1, 22.9, 22.7, 23.6, 23.8, 22.3, 21.8, 21.2, 20.0, 18.7, 17.7, 16.3, 15.2, 15.5, 15.2, 14.6, 12.0, 11.0, 12.8, 15.4, 18.8, 19.6, 21.3, 22.9, 23.8, 24.9, 26.2, 26.8, 26.3, 26.5, 26.3, 25.0, 21.8, 21.3, 16.6, 16.5, 16.1, 15.7, 14.1, 13.4, 13.1, 13.2, 13.2, 13.6, 14.8, 16.6, 17.4, 19.9, 20.4, 21.3, 21.7, 21.3, 22.4, 21.5, 21.5, 20.4, 18.0, 16.3, 15.7, 15.8, 15.2, 14.7, 14.4, 14.4, 14.7, 14.9, 14.5, 13.3, 13.2, 14.3, 16.2, 16.8, 18.2, 19.7, 19.3, 21.2, 14.4, 14.2, 13.9, 14.3, 14.1, 13.8, 13.9, 13.7, 13.8, 13.4, 13.1, 12.3, 12.9, 13.1, 13.3, 13.8, 13.5, 13.4, 14.1, 14.9, 15.5, 17.2, 17.8, 17.9, 19.1, 18.3, 18.0, 16.8, 14.7, 13.0, 12.2, 11.8, 10.9, 11.2, 9.8, 9.4, 8.5, 7.9, 9.1, 11.4, 12.1, 12.7, 13.4, 16.4, 18.5, 19.4, 21.0, 21.7, 22.5, 22.4, 21.8, 19.7, 18.4, 17.1, 17.0, 16.6, 15.4, 15.7, 16.4, 18.3, 16.5, 15.5, 13.8, 13.7, 14.6, 14.7, 15.2, 16.1, 16.4, 16.0, 17.0, 16.4, 18.8, 17.8, 18.0, 17.0, 16.4, 16.2, 14.5, 14.4, 14.9, 14.1, 13.9, 13.8, 12.4, 10.1, 10.8, 12.9, 14.3, 15.4, 17.7, 19.3, 19.9, 20.3, 21.2, 20.8, 21.6, 21.2, 21.3, 20.2, 18.2, 15.6, 13.9, 12.5, 12.3, 11.2, 10.6, 10.2, 9.9, 9.5, 10.5, 14.2, 16.7, 19.2, 21.4, 23.2, 24.5, 25.7, 25.9, 26.8, 26.3, 26.5, 26.2, 23.7, 20.8, 18.2, 16.0, 14.7, 13.7, 13.1, 12.0, 11.6, 10.8, 10.4, 12.3, 15.9, 18.0, 20.6, 22.8, 24.6, 26.0, 27.1, 27.5, 27.8, 28.2, 27.9, 27.7, 25.6, 22.2, 19.2, 17.8, 16.9, 15.6, 16.2, 15.5, 14.4, 14.0, 15.1, 15.6, 17.2, 19.1, 20.6, 21.5, 20.3, 20.5, 20.7, 20.1, 20.0, 20.1, 19.2, 18.1, 16.6, 16.0, 15.4, 15.2, 15.1, 14.9, 14.8, 13.6, 13.4, 13.2, 13.3, 13.3, 13.8, 14.9, 16.5, 17.1, 18.4, 19.0, 18.9, 19.1, 18.2, 18.8, 19.3, 18.7, 16.9, 14.5, 12.8, 12.3, 11.4, 10.7, 9.8, 9.7, 9.6, 9.0, 8.9, 9.6, 12.2, 14.5, 16.5, 16.6, 18.7, 19.4, 20.2, 21.7, 21.5, 21.4, 20.7, 21.1, 19.2, 17.1, 15.6, 14.6, 12.8, 10.9, 8.6, 6.7, 5.1, 4.8, 5.2, 5.1, 7.0, 10.8, 13.3, 14.7, 15.8, 17.2, 17.0, 16.7, 17.3, 15.6, 15.9, 15.8, 15.2, 14.3, 12.9, 10.7, 9.8, 9.5, 9.8, 9.0, 8.0, 7.5, 7.9, 8.1, 9.4, 11.8, 14.1, 15.9, 17.5, 18.1, 18.9, 19.9, 18.9, 18.7, 19.7, 19.3, 18.2, 16.3, 13.9, 11.5, 9.7, 10.2, 8.5, 8.2, 7.1, 5.9, 5.5, 6.4, 11.2, 14.2, 16.5, 18.0, 19.7, 21.1, 22.1, 21.9, 23.6, 23.7, 23.8, 22.3, 20.3, 18.6, 17.0, 15.4, 14.8, 13.6, 12.6, 11.4, 10.2, 9.8, 9.0, 9.9, 14.0, 17.1, 17.0, 19.9, 21.7, 23.3, 24.7, 25.2, 26.0, 26.4, 26.3, 25.2, 23.4, 22.0, 20.2, 19.3, 18.7, 18.3, 17.8, 17.4, 16.6, 16.3, 15.7, 15.2, 16.2, 18.7, 20.9, 22.4, 23.8, 25.2, 25.4, 26.1, 26.6, 27.2, 28.3, 27.4, 26.3, 23.9, 23.0, 23.7, 21.7, 19.7, 18.5, 18.2, 16.8, 16.1, 15.9, 15.9, 16.0, 17.0, 16.9, 17.5, 19.2, 19.6, 19.4, 20.1, 19.8, 19.6, 18.3, 18.4, 17.9, 16.9, 16.3, 15.7, 15.4, 15.0, 14.7, 14.5, 14.3, 14.4, 13.8, 13.9, 14.3, 15.0, 15.9, 17.8, 18.3, 18.4, 18.9, 19.0, 19.1, 19.5, 20.1, 19.7, 19.5, 17.8, 15.9, 15.4, 14.2, 13.2, 12.3, 11.3, 11.1, 10.4, 10.1, 11.1, 14.8, 17.7, 19.6, 21.6, 23.1, 24.3, 24.9, 25.3, 25.8, 26.3, 26.0, 24.6, 23.3, 22.9, 20.6, 19.2, 18.2, 17.5, 19.7, 18.0, 16.1, 15.3, 16.0, 15.5, 16.6, 17.4, 18.1, 17.3, 17.3, 17.4, 17.5, 18.5, 18.9, 19.0, 18.4, 18.8, 18.0, 16.8, 16.4, 16.0, 15.7, 15.4, 15.2, 15.0, 14.8, 14.6, 14.6, 14.9, 14.8, 14.7, 15.0, 15.7, 16.2, 16.5, 17.2, 18.2, 18.7, 19.0, 18.9, 17.7, 17.5, 16.6, 15.6, 15.0, 14.4, 14.2, 14.0, 14.0, 13.7, 13.7, 13.6, 13.5, 13.5, 13.7, 13.7, 13.8, 13.8, 14.2, 14.6, 14.8, 15.1, 14.7, 14.5, 14.5, 13.8, 13.8, 13.6, 13.6, 13.2, 12.6, 11.8, 11.2, 10.5, 10.4, 10.4, 10.0, 10.4, 11.4, 12.9, 13.9, 13.9, 14.2, 15.3, 15.0, 16.3, 17.3, 17.9, 16.7, 16.2, 14.6, 12.5, 11.1, 10.1, 9.5, 9.0, 8.7, 8.0, 8.5, 8.9, 10.5, 12.4, 13.7, 16.1, 17.5, 18.9, 20.5, 22.0, 21.8, 23.5, 22.5, 23.1, 21.7, 21.2, 20.8, 18.0, 16.3, 15.0, 14.4, 13.1, 12.3, 11.4, 10.7, 10.0, 11.7, 15.6, 17.8, 20.5, 22.7, 23.7, 25.2, 26.9, 27.5, 28.2, 28.3, 26.9, 26.8, 26.3, 24.8, 22.7, 21.4, 20.1, 18.6, 17.1, 15.9, 15.6, 14.5, 14.0, 15.2, 18.2, 20.7, 23.8, 25.5, 27.3, 28.1, 29.6, 30.4, 30.4, 31.1, 30.7, 30.0, 28.8, 27.0, 23.2, 23.7, 22.2, 20.7, 19.8, 19.2, 18.2, 18.7, 17.9, 17.3, 18.6, 19.8, 20.4, 21.6, 24.8, 26.3, 27.2, 24.5, 25.3, 23.7, 24.5, 25.0, 25.5, 25.0, 23.7, 20.8, 21.4, 21.3, 20.5, 20.2, 17.4, 16.8, 17.1, 16.8, 16.9, 18.4, 20.2, 22.0, 23.6, 23.8, 25.3, 23.3, 23.6, 25.1, 26.3, 24.8, 23.8, 21.3, 20.9, 20.0, 19.9, 19.4, 19.3, 18.4, 18.1, 17.2, 16.4, 15.5, 14.4, 14.9, 15.4, 15.2, 16.5, 17.1, 17.3, 18.8, 19.6, 19.8, 18.5, 18.4, 18.0, 17.6, 16.2, 15.7, 15.0, 15.8, 14.6, 14.2, 14.8, 13.0, 13.7, 13.3, 14.0, 14.8, 15.4, 16.8, 17.8, 18.5, 19.7, 19.7, 20.3, 20.5, 19.8, 20.7, 18.9, 18.7, 16.7, 13.9, 11.5, 10.6, 10.6, 10.3, 10.0, 9.5, 9.3, 10.8, 13.5, 16.5, 17.9, 19.7, 20.7, 21.6, 21.8, 22.7, 23.5, 23.7, 24.1, 23.7, 22.5, 20.3, 18.5, 17.6, 17.4, 16.4, 15.5, 15.3, 14.8, 14.0, 14.0, 15.4, 17.7, 19.6, 21.8, 23.7, 25.4, 27.5, 28.8, 29.5, 30.9, 30.8, 30.2, 29.6, 27.9, 26.7, 25.0, 23.2, 21.2, 19.5, 18.1, 17.2, 16.7, 16.4, 17.1, 16.5, 19.3, 21.2, 23.3, 24.8, 26.3, 27.6, 28.9, 28.5, 28.3, 28.6, 28.8, 26.5, 25.2, 23.5, 22.3, 20.2, 19.1, 18.2, 17.6, 16.8, 16.2, 16.1, 15.9, 16.8, 19.7, 21.5, 23.7, 25.7, 27.1, 28.5, 28.9, 30.5, 30.3, 28.3, 29.8, 29.8, 27.7, 25.4, 23.3, 21.7, 20.7, 19.8, 19.7, 19.2, 19.7, 19.6, 19.0, 19.4, 21.3, 23.2, 25.2, 26.5, 26.6, 28.2, 28.6, 29.2, 29.6, 29.6, 27.9, 25.1, 23.8, 22.6, 21.4, 20.0, 18.9, 17.6, 16.3, 15.0, 13.7, 12.6, 11.9, 12.0, 13.7, 14.9, 16.1, 16.7, 17.8, 19.0, 19.3, 20.4, 20.5, 21.2, 21.0, 20.0, 19.1, 18.1, 17.0, 15.1, 12.7, 11.2, 10.7, 9.8, 9.4, 9.2, 8.8, 10.0, 12.3, 15.1, 16.7, 17.9, 18.3, 18.8, 19.7, 20.1, 20.5, 20.6, 20.8, 20.2, 19.5, 18.2, 16.8, 16.0, 15.0, 13.3, 12.1, 11.2, 10.5, 9.9, 9.0, 10.2, 12.8, 15.4, 17.1, 18.6, 19.3, 20.7, 21.4, 21.9, 22.6, 23.4, 23.0, 22.6, 21.9, 20.7, 18.8, 17.7, 16.2, 15.3, 14.8, 13.6, 12.7, 11.8, 10.9, 11.6, 13.7, 16.6, 18.4, 19.6, 20.2, 21.4, 23.1, 21.9, 22.6, 22.3, 21.8, 22.7, 22.2, 21.2, 19.4, 17.8, 16.8, 15.4, 14.0, 12.7, 12.1, 11.7, 10.9, 12.1, 14.2, 17.2, 19.3, 21.1, 23.7, 24.7, 25.3, 25.5, 26.5, 27.3, 27.4, 26.6, 25.9, 24.2, 20.7, 18.1, 16.2, 15.0, 14.0, 13.2, 12.7, 12.2, 12.1, 13.7, 16.6, 18.4, 20.9, 23.5, 25.7, 27.0, 27.6, 28.3, 28.5, 28.1, 28.1, 26.6, 23.8, 23.0, 21.7, 19.9, 18.2, 16.7, 14.5, 13.8, 13.2, 12.9, 11.9, 12.3, 13.8, 14.6, 15.3, 16.4, 17.6, 18.7, 19.1, 19.8, 18.5, 19.3, 19.9, 19.5, 17.6, 16.7, 15.8, 15.1, 14.4, 13.2, 11.5, 11.6, 11.1, 10.4, 9.0, 10.2, 11.5, 13.7, 13.7, 13.1, 12.5, 12.8, 12.6, 12.7, 13.2, 15.2, 15.6, 16.6, 16.5, 16.0, 15.0, 14.3, 13.0, 12.7, 12.7, 12.7, 12.4, 11.9, 11.8, 11.5, 11.2, 11.2, 12.0, 12.6, 13.1, 13.9, 14.0, 14.4, 14.9, 14.9, 14.9, 15.6, 15.0, 13.9, 13.1, 12.6, 12.3, 12.1, 11.8, 11.6, 10.8, 10.3, 10.2, 10.1, 10.6, 11.3, 12.2, 13.3, 15.0, 14.7, 16.1, 16.7, 14.6, 16.2, 17.9, 16.5, 12.8, 12.0, 11.7, 11.5, 11.7, 11.3, 11.3, 11.1, 11.0, 10.9, 10.9, 10.8, 11.1, 11.7, 13.4, 14.3, 14.4, 15.6, 16.4, 16.3, 17.1, 16.5, 16.7, 16.4, 15.6, 15.0, 14.4, 13.8, 13.0, 12.6, 12.3, 12.0, 12.0, 11.8, 11.6, 11.2, 11.9, 12.7, 14.7, 14.7, 13.9, 15.0, 15.4, 15.3, 15.9, 15.9, 15.8, 15.5, 14.9, 14.5, 13.4, 11.1, 12.3, 11.8, 11.6, 11.3, 11.1, 10.7, 10.6, 10.9, 11.3, 12.0, 13.1, 14.9, 15.7, 15.7, 17.0, 18.3, 18.4, 18.2, 18.2, 18.6, 17.7, 16.3, 15.2, 14.2, 14.2, 14.7, 15.7, 16.7, 17.5, 17.8, 17.9, 18.1, 18.8, 19.7, 20.8, 23.0, 23.7, 23.9, 24.9, 25.6, 25.8, 25.4, 25.5, 25.4, 25.0, 24.0, 21.8, 19.0, 17.9, 17.4, 16.8, 18.6, 19.1, 18.9, 18.2, 17.5, 17.2, 17.4, 17.7, 19.6, 20.0, 20.6, 21.2, 22.4, 22.4, 23.6, 23.2, 22.3, 21.6, 21.0, 20.5, 19.7, 19.0, 18.5, 18.3, 16.8, 13.5, 12.3, 13.5, 14.3, 15.7, 17.3, 19.0, 20.7, 21.2, 20.5, 21.6, 22.0, 22.5, 22.5, 22.9, 22.5, 22.6, 21.1, 17.7, 16.0, 15.2, 14.3, 13.2, 13.1, 12.8, 13.7, 14.0, 15.0, 15.9, 17.7, 19.0, 20.1, 21.5, 23.2, 23.3, 23.2, 23.0, 22.4, 22.3, 22.0, 21.4, 20.4, 19.9, 19.3, 19.0, 17.3, 15.6, 16.5, 17.1, 17.2, 17.4, 17.5, 18.0, 17.1, 16.1, 15.4, 14.8, 14.9, 15.3, 16.7, 17.9, 18.8, 19.1, 19.1, 18.9, 18.4, 16.5, 14.8, 15.2, 14.0, 13.7, 13.1, 12.8, 12.6, 12.6, 12.8, 13.4, 15.3, 16.9, 19.2, 19.7, 20.3, 21.1, 22.0, 22.3, 22.7, 23.4, 22.7, 21.9, 20.5, 19.4, 18.8, 17.3, 16.6, 15.3, 14.8, 14.5, 13.8, 13.0, 13.5, 15.3, 17.4, 19.9, 20.7, 22.4, 22.7, 24.1, 25.6, 26.3, 25.4, 24.9, 23.9, 22.1, 20.2, 18.1, 16.6, 15.4, 14.7, 14.6, 14.0, 14.2, 14.4, 14.7, 14.6, 15.0, 15.6, 16.5, 16.7, 17.6, 19.5, 20.0, 20.3, 20.3, 21.1, 21.3, 21.0, 20.6, 20.3, 19.9, 18.6, 17.8, 18.5, 18.8, 18.9, 18.5, 18.1, 17.5, 17.1, 17.0, 17.5, 17.5, 17.9, 18.7, 19.6, 20.2, 19.7, 20.2, 20.6, 21.2, 21.4, 20.3, 19.7, 19.3, 18.9, 18.6, 18.3, 17.9, 17.5, 16.9, 16.5, 16.2, 16.3, 16.6, 16.7, 18.2, 18.5, 19.8, 21.0, 20.5, 21.1, 20.9, 20.3, 20.4, 20.9, 20.3, 19.3, 18.5, 17.7, 16.7, 15.4, 14.1, 12.7, 11.5, 11.1, 12.4, 12.4, 15.6, 16.9, 18.4, 19.8, 20.8, 22.1, 22.0, 21.6, 21.9, 22.9, 22.2, 21.9, 21.0, 20.1, 19.1, 18.3, 17.0, 16.1, 16.0, 14.1, 12.9, 12.5, 12.8, 15.5, 16.6, 18.9, 19.0, 20.2, 21.9, 22.5, 23.5, 23.8, 25.3, 24.7, 24.4, 23.2, 22.4, 20.3, 18.5, 18.3, 17.6, 17.6, 17.5, 17.5, 17.5, 16.6, 15.6, 15.4, 15.8, 16.3, 17.2, 17.6, 17.9, 18.6, 19.7, 20.9, 22.2, 21.2, 22.4, 21.5, 19.0, 17.4, 17.2, 15.8, 15.2, 13.4, 14.0, 14.0, 14.0, 13.3, 12.7, 13.0, 13.3, 14.1, 14.4, 13.3, 14.7, 15.5, 18.1, 19.0, 19.4, 18.0, 16.8, 14.1, 15.0, 14.1, 12.8, 13.0, 13.1, 13.2, 12.4, 11.8, 11.8, 11.7, 10.6, 10.8, 13.1, 13.6, 16.0, 17.4, 18.4, 20.1, 19.3, 19.4, 20.9, 22.5, 20.8, 18.3, 18.0, 16.0, 15.3, 15.8, 15.5, 15.2, 15.3, 15.1, 14.6, 13.9, 14.0, 13.7, 15.0, 16.4, 16.7, 17.7, 18.7, 19.7, 19.9, 20.7, 22.2, 22.6, 22.4, 22.1, 22.4, 21.3, 20.9, 19.6, 17.0, 16.4, 16.1, 16.1, 16.8, 16.4, 16.8, 16.5, 17.1, 19.2, 19.4, 20.7, 22.4, 24.0, 24.1, 24.8, 26.0, 26.9, 27.3, 27.1, 26.6, 23.9, 21.4, 19.2, 18.7, 16.9, 16.6, 16.2, 15.2, 14.7, 15.2, 18.1, 21.1, 23.1, 24.9, 26.4, 28.1, 29.6, 30.9, 31.1, 31.7, 31.9, 32.0, 31.3, 29.8, 27.4, 23.3, 22.0, 20.4, 19.0, 18.9, 18.6, 17.5, 17.2, 17.1, 18.6, 22.7, 24.5, 27.7, 29.1, 32.0, 33.4, 34.1, 35.7, 35.7, 36.3, 35.8, 35.7, 34.0, 28.3, 24.9, 22.8, 21.1, 20.2, 19.9, 19.1, 18.4, 18.0, 17.3, 20.3, 24.9, 27.4, 28.6, 29.5, 30.8, 32.3, 33.4, 34.1, 34.0, 34.9, 34.7, 34.2, 31.9, 27.9, 30.0, 27.2, 25.7, 24.5, 25.7, 25.9, 24.4, 23.2, 22.0, 21.5, 22.2, 22.2, 20.7, 23.1, 24.8, 23.6, 26.0, 26.7, 27.6, 26.4, 27.0, 26.8, 26.4, 24.9, 23.2, 21.8, 20.0, 20.5, 19.9, 19.3, 19.6, 18.9, 18.8, 18.8, 19.8, 20.5, 21.3, 22.1, 24.4, 25.5, 26.8, 27.1, 26.9, 28.7, 28.7, 28.4, 27.8, 27.2, 24.9, 23.5, 22.0, 21.0, 20.3, 19.6, 19.0, 18.6, 18.0, 18.7, 17.8, 17.2, 20.4, 20.5, 18.6, 17.5, 21.8, 24.1, 23.7, 23.3, 23.3, 24.3, 23.7, 21.9, 20.5, 19.7, 19.4, 18.9, 18.8, 18.4, 18.0, 17.7, 17.5, 17.5, 20.1, 21.8, 24.4, 27.0, 28.4, 28.2, 24.8, 24.7, 25.3, 25.0, 26.9, 25.4, 25.9, 23.7, 22.1, 21.3, 21.1, 20.8, 20.7, 19.5, 17.8, 18.3, 18.2, 18.6, 19.0, 18.4, 19.2, 19.6, 19.6, 20.9, 21.7, 22.0, 21.0, 19.9, 18.4, 17.8, 16.2, 16.1, 16.0, 15.8, 15.8, 15.8, 15.9, 15.8, 15.6, 15.3, 15.2, 15.6, 16.3, 17.0, 18.0, 20.7, 19.9, 21.4, 23.2, 23.5, 23.8, 22.6, 24.3, 23.2, 22.6, 20.8, 16.7, 15.4, 14.7, 13.2, 13.5, 12.3, 11.7, 11.6, 12.6, 13.9, 17.1, 17.3, 17.1, 20.3, 22.2, 23.4, 25.1, 25.9, 24.0, 22.5, 21.7, 19.4, 17.4, 17.8, 17.5, 17.5, 18.0, 18.5, 19.0, 19.6, 20.1, 20.2, 20.3, 20.2, 21.1, 22.5, 24.7, 25.7, 27.9, 29.3, 30.7, 30.1, 22.4, 25.3, 26.8, 26.6, 22.7, 20.7, 20.3, 19.6, 19.4, 19.2, 19.0, 19.1, 19.4, 19.5, 19.5, 19.5, 19.8, 20.3, 21.4, 22.1, 22.9, 23.7, 24.4, 25.7, 25.1, 25.6, 25.9, 25.2, 24.5, 23.0, 20.9, 19.6, 18.0, 16.7, 15.7, 15.7, 14.7, 12.8, 12.1, 12.9, 15.6, 17.8, 19.8, 21.2, 22.9, 23.9, 24.4, 26.0, 26.3, 26.2, 25.7, 24.0, 23.0, 21.7, 20.2, 18.5, 17.6, 17.1, 16.6, 16.4, 16.2, 14.9, 14.7, 14.8, 15.5, 16.7, 17.0, 17.7, 18.4, 18.8, 19.3, 21.0, 21.1, 16.5, 17.7, 18.1, 18.1, 17.0, 17.0, 16.7, 15.4, 13.9, 12.8, 11.9, 12.1, 11.8, 11.4, 11.8, 14.0, 15.6, 17.2, 18.4, 19.8, 20.2, 22.1, 22.0, 21.7, 22.5, 22.2, 22.1, 21.3, 20.2, 18.4, 17.5, 16.2, 15.2, 14.4, 13.4, 12.7, 12.0, 11.4, 11.8, 14.3, 17.7, 19.6, 21.1, 22.0, 22.9, 23.9, 24.3, 25.0, 25.7, 25.4, 24.9, 24.0, 22.2, 21.0, 19.7, 17.3, 16.7, 18.9, 18.7, 18.6, 18.0, 16.0, 15.9, 18.9, 20.8, 22.4, 24.1, 24.8, 24.9, 25.9, 26.3, 27.7, 27.8, 27.2, 27.0, 25.9, 23.8, 20.8, 19.5, 17.9, 16.8, 15.6, 14.9, 14.0, 14.2, 12.9, 14.3, 17.3, 20.0, 22.4, 24.4, 25.8, 28.1, 28.1, 29.0, 29.9, 29.6, 29.8, 29.2, 28.2, 25.5, 22.1, 20.0, 18.8, 17.8, 16.8, 16.0, 15.4, 14.9, 14.6, 14.6, 18.0, 19.9, 22.7, 24.4, 26.5, 28.5, 29.2, 30.6, 31.5, 30.4, 30.1, 29.8, 29.0, 27.0, 24.6, 24.7, 23.9, 23.1, 22.3, 21.6, 20.8, 20.5, 19.7, 19.4, 20.0, 22.5, 24.1, 25.7, 26.6, 27.9, 27.7, 28.2, 28.3, 29.2, 28.4, 28.3, 26.8, 25.6, 24.1, 22.5, 21.8, 21.6, 22.2, 23.1, 23.8, 24.0, 23.8, 23.8, 23.9, 24.0, 24.3, 23.8, 24.0, 25.1, 25.6, 21.5, 21.9, 23.0, 22.9, 22.6, 22.6, 21.2, 19.4, 18.6, 19.2, 18.7, 18.6, 18.8, 18.6, 18.3, 18.1, 17.5, 18.0, 19.0, 20.1, 21.5, 20.4, 19.7, 19.6, 21.0, 21.9, 22.9, 23.6, 22.8, 21.7, 20.7, 18.6, 17.6, 17.1, 18.1, 17.2, 15.8, 15.4, 15.0, 15.3, 15.4, 16.4, 18.7, 19.8, 20.2, 20.9, 21.8, 21.9, 23.0, 22.5, 21.0, 22.3, 21.2, 20.7, 19.6, 18.0, 17.3, 16.0, 15.2, 15.8, 15.8, 16.0, 16.0, 16.1, 15.9, 16.5, 17.2, 17.5, 17.9, 20.7, 22.1, 21.4, 22.1, 21.1, 21.6, 21.6, 20.7, 19.7, 19.0, 18.4, 18.4, 18.2, 18.2, 18.1, 18.0, 17.8, 17.6, 17.3, 17.1, 17.3, 17.4, 17.8, 18.0, 18.7, 20.5, 20.7, 19.9, 19.5, 19.0, 19.2, 19.5, 19.4, 18.5, 17.9, 17.9, 17.6, 18.1, 18.5, 19.0, 18.0, 17.5, 18.0, 17.7, 18.0, 19.0, 19.3, 20.8, 21.8, 21.8, 22.3, 23.2, 22.7, 23.4, 24.3, 22.5, 18.6, 17.8, 17.0, 16.2, 16.5, 16.6, 16.3, 15.9, 16.3, 16.7, 16.4, 16.5, 16.5, 17.4, 18.7, 20.2, 20.7, 22.2, 23.9, 22.7, 21.4, 21.3, 21.0, 20.7, 19.2, 18.3, 17.2, 17.2, 17.2, 16.7, 15.9, 15.8, 15.7, 15.0, 15.7, 14.7, 15.9, 16.8, 17.7, 17.1, 17.3, 18.3, 17.6, 20.2, 20.1, 20.8, 19.6, 17.5, 14.9, 13.8, 14.2, 14.0, 13.6, 13.0, 13.0, 13.0, 12.3, 11.1, 10.8, 10.2, 12.5, 14.5, 15.4, 16.6, 17.7, 18.9, 20.8, 21.1, 21.7, 22.5, 20.8, 21.0, 19.5, 17.4, 15.0, 13.7, 12.6, 11.6, 11.1, 10.3, 10.0, 9.6, 9.4, 9.2, 12.4, 14.8, 17.9, 19.7, 21.8, 22.1, 22.4, 23.8, 24.3, 25.0, 25.1, 24.0, 23.3, 21.1, 19.3, 18.3, 17.3, 16.5, 15.9, 15.6, 15.0, 16.0, 15.8, 15.5, 15.9, 17.5, 18.8, 20.9, 23.8, 24.7, 26.8, 26.8, 28.0, 28.6, 28.9, 28.3, 26.9, 25.1, 22.2, 20.3, 19.1, 18.4, 17.4, 16.7, 16.5, 15.9, 15.1, 15.6, 18.7, 21.0, 23.3, 25.3, 28.6, 29.7, 30.5, 31.9, 32.0, 32.9, 32.5, 32.3, 31.0, 28.4, 26.1, 25.4, 22.5, 20.8, 20.0, 19.2, 18.7, 18.4, 18.4, 17.9, 21.0, 24.2, 26.4, 27.8, 30.3, 31.6, 32.8, 33.7, 34.6, 34.2, 34.8, 34.2, 30.9, 27.4, 24.3, 22.4, 22.2, 22.0, 20.6, 19.4, 19.9, 18.8, 18.8, 19.2, 21.6, 23.8, 26.2, 27.2, 29.1, 30.0, 29.6, 29.9, 28.5, 27.8, 26.3, 26.0, 25.2, 24.6, 23.0, 21.8, 21.1, 20.5, 19.8, 18.9, 19.2, 19.2, 19.0, 18.9, 19.2, 20.7, 22.1, 23.6, 24.9, 26.1, 26.0, 26.9, 27.1, 27.1, 26.3, 24.8, 23.5, 21.6, 19.7, 18.9, 18.8, 18.6, 19.2, 19.2, 18.9, 18.2, 18.2, 18.1, 20.7, 22.9, 23.6, 24.6, 24.5, 25.0, 25.5, 25.8, 27.5, 28.3, 28.2, 28.1, 26.9, 25.2, 23.6, 22.1, 20.2, 18.5, 17.0, 15.9, 14.9, 14.5, 14.4, 13.5, 14.6, 17.9, 20.9, 22.1, 23.8, 24.3, 24.6, 25.2, 25.9, 25.8, 25.1, 24.5, 24.0, 22.8, 21.3, 19.9, 18.2, 18.9, 18.9, 18.2, 17.4, 17.0, 16.2, 15.9, 17.2, 20.8, 23.0, 24.8, 25.7, 26.9, 27.7, 28.5, 29.0, 29.3, 28.9, 28.2, 26.9, 24.4, 21.0, 20.2, 19.3, 19.4, 17.3, 17.6, 17.9, 18.2, 17.3, 16.4, 17.8, 20.7, 22.7, 24.0, 25.3, 25.7, 27.5, 27.8, 29.0, 29.6, 29.3, 28.3, 26.4, 23.1, 21.3, 20.9, 22.4, 21.2, 19.6, 18.4, 17.7, 17.5, 17.9, 18.0, 18.3, 18.9, 20.0, 21.0, 20.9, 20.9, 21.8, 24.9, 24.8, 24.4, 24.6, 24.5, 21.9, 21.7, 20.4, 19.8, 19.4, 18.9, 18.3, 18.0, 17.4, 16.8, 16.5, 16.8, 17.5, 17.9, 18.7, 19.8, 21.4, 22.9, 23.8, 25.0, 25.0, 25.4, 24.8, 24.6, 24.1, 23.4, 21.9, 20.1, 19.3, 18.5, 17.7, 17.8, 17.9, 17.4, 16.5, 16.9, 17.5, 17.6, 18.3, 19.6, 21.1, 22.2, 22.6, 24.2, 25.3, 25.9, 26.2, 25.8, 24.2, 21.2, 19.4, 18.7, 18.8, 19.4, 21.2, 19.8, 18.7, 17.8, 16.5, 15.7, 16.0, 16.7, 16.9, 17.7, 19.9, 21.7, 23.1, 24.1, 22.6, 23.1, 23.3, 22.2, 21.7, 19.7, 19.3, 18.2, 17.1, 16.4, 16.6, 16.0, 15.8, 14.8, 13.6, 12.9, 13.9, 16.9, 19.4, 21.4, 22.2, 22.6, 22.0, 22.5, 24.1, 23.5, 22.6, 22.9, 21.5, 20.0, 17.8, 15.4, 14.9, 13.8, 13.8, 13.9, 13.4, 12.6, 12.7, 13.4, 14.6, 16.0, 17.2, 19.5, 22.0, 23.7, 24.1, 20.7, 20.2, 22.1, 21.7, 21.9, 21.1, 19.4, 18.7, 17.6, 17.4, 16.7, 15.3, 14.2, 13.4, 13.8, 13.8, 13.8, 14.3, 15.7, 16.2, 17.6, 20.2, 21.9, 23.3, 23.4, 23.1, 23.0, 22.9, 22.3, 21.2, 20.1, 19.1, 18.3, 17.0, 15.8, 15.5, 15.3, 15.2, 15.0, 14.9, 15.0, 15.1, 15.3, 15.0, 14.9, 15.1, 16.2, 19.0, 19.2, 18.6, 18.3, 18.7, 18.5, 17.1, 15.6, 13.6, 11.9, 12.1, 13.3, 12.4, 11.9, 12.3, 12.4, 12.5, 11.9, 12.2, 13.5, 15.3, 16.9, 18.3, 19.2, 19.2, 21.1, 19.7, 19.1, 19.3, 18.6, 17.9, 17.0, 16.2, 15.2, 14.7, 14.3, 13.8, 12.8, 12.6, 12.2, 12.0, 12.0, 12.2, 12.8, 13.5, 14.7, 14.4, 15.1, 15.8, 15.9, 16.3, 17.2, 17.1, 17.2, 16.7, 15.9, 15.3, 14.8, 14.7, 14.9, 15.2, 15.4, 15.4, 15.1, 15.1, 14.6, 14.7, 15.0, 15.6, 16.3, 17.4, 17.8, 18.6, 19.3, 21.2, 22.0, 22.2, 22.7, 21.7, 20.5, 18.9, 17.6, 16.4, 15.6, 14.5, 14.3, 14.4, 14.5, 15.2, 15.4, 15.6, 16.3, 17.0, 18.6, 19.4, 21.8, 23.7, 23.6, 22.5, 21.4, 20.8, 17.3, 15.8, 16.0, 16.0, 16.2, 15.3, 14.7, 13.6, 13.3, 13.0, 13.3, 12.8, 12.6, 13.6, 14.7, 15.5, 15.6, 16.9, 15.5, 14.9, 15.2, 15.7, 16.7, 15.7, 15.1, 14.5, 14.2, 14.0, 13.8, 13.5, 13.8, 13.2, 13.1, 13.1, 12.9, 12.8, 13.1, 13.3, 14.1, 15.0, 15.6, 16.1, 16.7, 18.0, 17.5, 17.8, 18.9, 16.8, 16.3, 15.9, 15.6, 14.3, 14.2, 12.6, 12.0, 12.3, 12.4, 12.1, 12.1, 12.1, 12.0, 12.0, 12.4, 14.1, 15.0, 16.3, 17.0, 18.3, 18.8, 16.4, 16.3, 16.1, 15.8, 14.9, 14.6, 14.6, 13.5, 13.1, 12.7, 12.6, 12.3, 12.5, 12.4, 11.4, 10.8, 11.2, 12.1, 14.8, 14.5, 14.6, 15.1, 16.8, 18.0, 17.8, 16.5, 17.4, 17.0, 16.2, 14.8, 13.7, 12.5, 11.1, 10.7, 10.5, 10.1, 10.4, 10.7, 10.3, 10.3, 10.6, 12.1, 12.9, 14.3, 14.5, 14.7, 15.5, 16.2, 15.4, 14.8, 14.8, 14.0, 13.8, 13.6, 13.6, 14.2, 14.4, 14.4, 14.3, 13.4, 11.8, 13.0, 12.6, 12.9, 12.5, 12.8, 14.6, 14.8, 16.9, 16.4, 16.6, 16.8, 16.8, 16.9, 16.0, 16.0, 15.4, 14.9, 14.5, 13.3, 12.2, 11.4, 10.8, 11.2, 11.2, 11.0, 10.8, 10.9, 11.6, 13.1, 14.5, 15.9, 18.5, 19.0, 20.6, 21.5, 21.7, 22.4, 22.4, 21.6, 19.7, 17.2, 15.3, 14.3, 13.5, 12.6, 12.3, 12.0, 11.3, 11.0, 10.7, 10.1, 10.1, 13.3, 15.9, 18.6, 20.8, 22.1, 22.9, 23.7, 24.3, 24.4, 24.6, 23.1, 22.3, 19.7, 18.2, 17.3, 16.6, 15.8, 15.4, 14.8, 14.2, 13.8, 13.2, 12.8, 12.8, 15.1, 16.8, 19.1, 22.2, 23.7, 25.6, 26.3, 26.1, 27.0, 26.5, 25.4, 23.6, 21.9, 20.3, 18.9, 17.9, 17.1, 16.4, 15.7, 15.4, 15.0, 14.5, 13.4, 12.9, 16.1, 18.6, 21.0, 23.1, 24.6, 25.0, 26.5, 27.3, 26.9, 26.7, 26.0, 23.3, 20.8, 18.7, 17.4, 16.4, 15.6, 15.6, 14.8, 14.3, 13.6, 13.8, 13.0, 12.6, 16.4, 19.0, 21.0, 23.9, 25.9, 26.3, 27.3, 27.3, 27.1, 26.4, 25.6, 23.4, 21.0, 19.5, 18.1, 17.2, 17.1, 16.9, 16.5, 17.2, 18.9, 17.3, 16.7, 16.5, 16.7, 17.6, 19.4, 20.0, 20.0, 20.2, 21.6, 22.5, 23.2, 21.9, 20.9, 19.2, 17.7, 16.3, 15.3, 14.5, 14.5, 14.7, 14.4, 14.2, 13.3, 12.3, 11.8, 11.8, 13.0, 15.1, 16.2, 16.8, 17.9, 20.3, 22.0, 21.7, 21.5, 21.6, 20.8, 20.4, 19.2, 18.0, 16.9, 16.0, 15.2, 15.4, 15.2, 14.8, 14.8, 14.2, 13.4, 13.5, 14.5, 16.2, 18.5, 20.5, 22.1, 23.5, 24.3, 24.6, 25.2, 24.7, 23.8, 22.3, 20.3, 18.8, 17.9, 17.7, 17.5, 17.6, 19.6, 17.8, 16.9, 17.3, 14.6, 13.9, 14.0, 14.0, 14.8, 15.0, 14.8, 16.0, 16.8, 18.1, 16.8, 16.2, 14.7, 14.4, 13.5, 13.5, 13.4, 13.6, 14.2, 14.5, 14.7, 14.7, 14.6, 14.3, 14.1, 13.9, 13.8, 14.0, 14.4, 14.6, 15.0, 15.5, 16.4, 16.6, 16.1, 15.6, 15.6, 15.3, 15.0, 15.0, 14.7, 14.8, 14.6, 14.5, 14.3, 14.4, 14.3, 14.4, 14.3, 14.0, 13.9, 14.9, 16.8, 16.8, 16.9, 17.1, 16.9, 18.4, 18.4, 18.7, 18.1, 17.0, 15.8, 14.8, 14.7, 13.7, 12.8, 12.0, 11.4, 10.6, 10.3, 9.8, 9.7, 9.7, 11.7, 14.6, 16.9, 19.3, 21.5, 22.8, 23.4, 22.8, 21.9, 20.6, 19.1, 17.1, 15.4, 16.1, 15.4, 13.7, 14.1, 13.8, 13.1, 13.0, 13.1, 12.5, 12.1, 12.3, 13.3, 14.1, 14.5, 16.8, 18.4, 17.9, 18.0, 17.3, 17.2, 17.0, 16.9, 16.3, 15.9, 15.8, 14.8, 14.5, 14.5, 14.4, 14.4, 13.9, 13.5, 13.4, 13.0, 12.8, 12.4, 12.3, 12.6, 13.1, 13.5, 13.7, 14.2, 14.5, 14.3, 14.0, 14.0, 13.8, 13.5, 13.2, 12.6, 12.1, 11.8, 11.7, 11.6, 11.5, 11.6, 11.6, 11.6, 11.6, 11.6, 13.1, 14.6, 15.5, 17.4, 18.2, 18.7, 19.1, 18.9, 18.3, 18.0, 16.7, 15.3, 14.9, 13.1, 12.9, 12.3, 11.2, 11.8, 11.5, 10.9, 10.1, 9.9, 10.6, 11.6, 13.5, 15.3, 16.6, 16.5, 17.2, 18.3, 18.3, 17.9, 17.4, 16.9, 15.4, 14.6, 12.6, 12.3, 12.9, 12.3, 10.2, 9.8, 8.5, 8.1, 8.3, 8.0, 7.4, 9.7, 13.7, 15.5, 16.4, 17.7, 18.8, 19.9, 21.0, 21.0, 21.4, 20.4, 17.1, 15.4, 13.5, 12.2, 11.8, 11.5, 11.1, 10.7, 10.8, 11.4, 11.6, 11.0, 12.0, 12.6, 13.1, 13.9, 15.3, 16.4, 16.5, 18.0, 18.5, 17.9, 18.0, 17.7, 16.2, 15.0, 13.9, 13.1, 12.4, 11.8, 11.4, 11.0, 10.5, 10.1, 9.9, 9.0, 9.2, 9.4, 9.7, 10.1, 10.3, 10.7, 13.0, 15.0, 13.8, 13.3, 13.3, 12.9, 12.1, 11.8, 11.5, 11.3, 11.2, 11.1, 10.9, 11.1, 11.2, 11.1, 10.8, 10.9, 11.2, 11.7, 12.2, 12.5, 13.8, 15.7, 16.2, 15.5, 15.4, 15.2, 14.5, 13.9, 13.8, 13.9, 13.6, 13.7, 13.3, 12.8, 12.8, 12.5, 12.6, 12.7, 12.5, 12.3, 12.6, 12.9, 15.5, 16.4, 17.6, 18.3, 18.9, 18.3, 18.6, 18.4, 17.8, 17.2, 16.6, 15.0, 13.8, 13.7, 12.6, 12.5, 12.8, 13.3, 14.0, 14.2, 14.2, 14.2, 14.0, 14.5, 15.0, 15.1, 16.6, 16.8, 17.5, 18.1, 18.6, 16.4, 18.2, 17.0, 16.0, 15.7, 13.8, 13.3, 12.7, 11.8, 11.0, 10.9, 10.5, 10.4, 10.2, 10.2, 10.0, 11.5, 13.0, 14.3, 15.7, 17.1, 18.3, 17.1, 17.8, 16.9, 16.4, 15.6, 14.8, 14.2, 14.2, 13.4, 12.1, 12.3, 12.4, 12.6, 12.6, 11.7, 11.2, 11.4, 11.8, 12.1, 13.1, 14.2, 14.9, 15.0, 15.1, 14.8, 15.2, 15.7, 15.9, 14.6, 12.9, 12.1, 12.0, 11.7, 12.1, 12.2, 11.8, 11.9, 11.3, 13.4, 12.3, 12.2, 11.1, 12.3, 12.9, 14.4, 16.7, 17.6, 19.3, 19.2, 18.4, 19.0, 17.9, 16.2, 14.5, 13.4, 12.7, 12.3, 12.0, 11.5, 10.5, 10.1, 10.0, 10.0, 9.1, 8.9, 8.7, 10.3, 13.5, 15.2, 17.2, 18.4, 19.3, 19.7, 18.9, 19.2, 18.5, 15.9, 13.7, 12.4, 11.3, 10.0, 9.7, 10.1, 9.6, 9.9, 9.2, 8.9, 8.0, 7.3, 7.6, 10.1, 15.0, 16.8, 17.8, 20.2, 21.8, 23.0, 23.0, 22.7, 22.1, 20.0, 17.9, 16.1, 15.4, 16.0, 15.4, 15.0, 16.0, 15.4, 14.6, 15.4, 15.2, 15.2, 14.6, 16.1, 16.9, 20.5, 22.9, 24.5, 25.8, 26.5, 26.6, 26.3, 24.5, 21.1, 19.0, 18.5, 17.8, 17.3, 15.8, 13.5, 10.8, 8.3, 6.2, 5.5, 5.7, 5.3, 5.1, 5.7, 7.3, 9.8, 11.9, 13.5, 14.6, 15.1, 16.0, 15.7, 14.5, 13.3, 10.9, 9.6, 8.8, 7.3, 7.0, 7.9, 7.9, 7.8, 8.1, 7.9, 7.6, 7.0, 7.3, 7.5, 7.9, 8.6, 9.7, 10.6, 11.3, 12.5, 12.8, 12.2, 11.5, 10.9, 10.9, 10.9, 11.0, 11.2, 11.2, 11.5, 11.7, 11.8, 12.0, 12.1, 11.9, 11.9, 11.8, 12.0, 12.7, 13.3, 14.4, 15.2, 14.6, 14.6, 15.5, 15.4, 14.9, 14.5, 13.9, 13.8, 13.3, 13.2, 13.3, 13.2, 13.3, 13.5, 13.3, 13.1, 13.1, 13.0, 13.0, 13.1, 13.3, 13.8, 14.2, 13.8, 14.4, 15.0, 15.2, 15.2, 14.9, 14.6, 13.8, 13.5, 13.8, 13.5, 13.3, 13.1, 13.1, 12.6, 12.5, 12.2, 12.1, 12.0, 11.9, 12.0, 12.8, 13.8, 15.6, 15.6, 16.6, 16.9, 16.6, 16.4, 16.7, 15.8, 13.9, 12.9, 12.6, 12.2, 12.7, 13.1, 13.3, 13.2, 13.4, 13.4, 13.0, 12.5, 12.2, 11.9, 12.1, 12.7, 13.1, 14.0, 14.1, 15.0, 15.3, 15.6, 15.3, 13.7, 11.8, 10.3, 8.4, 9.0, 7.3, 6.8, 6.4, 6.1, 5.9, 7.0, 7.4, 7.0, 5.7, 5.4, 7.8, 9.4, 10.9, 12.9, 14.7, 16.1, 15.9, 16.3, 15.6, 13.7, 11.5, 10.1, 8.7, 8.0, 6.9, 6.6, 7.5, 7.3, 6.1, 5.2, 4.4, 4.3, 4.0, 4.2, 5.8, 7.8, 10.5, 13.1, 14.3, 16.0, 15.3, 15.2, 15.0, 13.0, 12.8, 10.9, 9.7, 8.7, 7.7, 7.1, 6.6, 6.2, 6.0, 4.8, 3.7, 3.4, 3.2, 3.3, 5.7, 9.0, 12.3, 14.2, 16.1, 15.8, 15.8, 15.7, 14.5, 14.3, 12.6, 11.6, 10.5, 10.3, 10.0, 9.5, 9.0, 7.1, 7.4, 6.8, 5.7, 4.6, 3.7, 3.4, 7.2, 9.3, 11.4, 13.1, 14.4, 14.6, 15.2, 14.5, 13.5, 11.0, 9.8, 7.1, 4.9, 5.1, 7.0, 6.1, 5.8, 4.7, 5.6, 5.6, 4.6, 4.4, 2.8, 2.2, 7.1, 9.5, 10.6, 11.2, 12.4, 12.4, 12.6, 12.2, 11.3, 9.5, 8.4, 7.3, 6.1, 5.7, 5.4, 4.8, 5.3, 4.2, 2.5, 1.8, 1.6, 1.3, 0.7, 1.4, 5.7, 7.8, 9.1, 9.8, 10.7, 11.2, 11.4, 11.4, 10.6, 8.9, 8.4, 8.0, 7.1, 6.6, 5.9, 5.4, 4.7, 4.0, 3.6, 3.5, 3.0, 2.6, 1.4, 2.5, 5.0, 6.9, 8.7, 9.3, 10.4, 11.2, 10.8, 10.8, 9.8, 8.6, 7.3, 7.0, 5.8, 6.2, 6.7, 6.5, 6.7, 6.3, 5.7, 4.7, 4.7, 5.3, 5.6, 5.3, 5.3, 6.1, 7.5, 8.3, 9.9, 10.9, 10.9, 11.1, 9.9, 9.0, 9.2, 9.2, 8.7, 8.8, 8.6, 8.3, 8.2, 8.5, 7.8, 6.7, 7.1, 6.6, 6.5, 6.7, 7.7, 8.7, 10.3, 10.4, 10.6, 11.6, 11.9, 12.7, 11.9, 11.0, 9.9, 9.6, 8.9, 8.6, 8.2, 7.7, 6.4, 5.4, 4.2, 3.6, 3.7, 2.8, 2.9, 3.8, 6.1, 8.3, 8.8, 11.5, 14.1, 16.0, 15.8, 15.4, 14.8, 13.8, 10.9, 11.1, 11.4, 9.6, 9.8, 10.7, 9.6, 10.4, 9.5, 9.3, 10.0, 10.0, 10.4, 11.3, 12.2, 13.1, 13.7, 13.7, 14.2, 14.5, 15.0, 15.8, 14.4, 11.7, 10.7, 9.3, 9.5, 9.8, 9.0, 7.9, 8.3, 7.7, 7.2, 7.2, 6.0, 4.4, 4.1, 5.0, 8.6, 13.7, 14.5, 14.1, 13.9, 13.3, 13.1, 12.0, 11.7, 11.1, 11.1, 11.4, 11.1, 10.8, 11.1, 11.2, 11.0, 10.9, 10.8, 10.2, 10.1, 10.5, 10.1, 10.2, 10.7, 11.2, 11.3, 11.4, 12.2, 12.5, 12.8, 12.5, 12.3, 11.5, 10.5, 10.3, 10.1, 10.2, 9.3, 9.3, 8.9, 8.8, 7.7, 8.1, 7.6, 8.3, 7.0, 7.0, 9.2, 12.2, 14.4, 16.4, 17.2, 17.2, 17.1, 16.7, 16.0, 15.4, 14.8, 15.1, 13.8, 13.3, 10.3, 8.8, 7.7, 7.1, 7.4, 6.5, 7.1, 6.6, 6.6, 6.8, 8.7, 10.9, 13.3, 14.8, 15.7, 15.8, 16.5, 17.0, 15.7, 12.9, 10.1, 8.9, 7.5, 6.6, 5.4, 5.1, 4.5, 3.7, 2.7, 2.7, 2.4, 1.6, 2.7, 3.2, 4.9, 5.2, 7.0, 8.3, 11.9, 13.5, 13.2, 13.3, 13.3, 11.9, 10.6, 10.1, 10.3, 9.7, 8.5, 8.4, 8.7, 8.9, 8.8, 8.7, 8.6, 7.8, 7.0, 6.7, 6.9, 7.7, 9.7, 10.9, 12.5, 14.9, 15.8, 16.3, 14.9, 12.4, 10.7, 9.4, 8.5, 8.2, 9.1, 10.3, 11.8, 12.9, 13.6, 13.4, 13.2, 12.8, 12.3, 11.7, 11.6, 11.8, 12.3, 13.4, 13.8, 14.1, 14.4, 14.4, 13.6, 12.9, 11.6, 11.5, 11.9, 11.5, 10.3, 9.8, 8.7, 7.9, 7.0, 6.6, 6.4, 7.1, 7.6, 7.8, 8.2, 9.5, 12.2, 12.3, 13.1, 13.6, 14.3, 13.7, 11.7, 10.0, 7.5, 6.1, 5.0, 5.0, 4.2, 4.2, 3.7, 4.2, 3.2, 3.3, 3.0, 3.2, 4.5, 5.4, 6.3, 7.0, 7.3, 7.8, 8.5, 8.9, 9.2, 9.7, 9.3, 9.2, 9.0, 9.1, 8.1, 7.9, 7.4, 7.2, 7.4, 7.4, 6.7, 6.0, 6.2, 5.6, 5.1, 5.4, 5.8, 6.9, 8.6, 9.3, 8.7, 8.8, 9.3, 8.8, 8.2, 6.9, 5.7, 5.8, 6.7, 7.1, 8.0, 8.3, 8.6, 8.6, 9.1, 9.1, 9.3, 9.2, 9.0, 8.9, 9.2, 9.3, 8.9, 8.3, 9.6, 8.8, 9.5, 8.4, 8.0, 7.8, 5.9, 5.8, 4.9, 4.5, 3.4, 2.5, 1.6, 1.2, 1.2, 1.2, 1.7, 1.7, 1.7, 1.7, 1.5, 2.3, 2.6, 3.8, 4.1, 4.2, 4.8, 4.4, 3.5, 2.0, 0.8, -0.3, -0.9, -1.2, -1.7, -2.8, -3.2, -3.1, -3.5, -3.4, -3.8, -4.1, -4.1, -4.3, -2.9, 0.5, 2.5, 4.0, 4.4, 4.7, 4.0, 3.9, 2.5, 1.1, -0.5, -1.2, -2.0, -3.0, -4.0, -4.4, -4.4, -5.2, -4.7, -5.2, -6.1, -6.6, -6.5, -5.0, -3.5, -2.1, -0.9, 0.8, 2.4, 3.5, 4.0, 3.8, 2.6, 0.3, -1.0, -1.4, -1.7, -1.4, -1.8, -1.9, -1.9, -2.1, -2.3, -2.5, -3.0, -1.9, -1.2, -0.8, 0.0, 0.8, 1.1, 1.5, 2.1, 2.2, 2.4, 2.5, 2.6, 2.6, 2.7, 3.0, 3.0, 3.0, 2.8, 2.9, 3.0, 3.1, 3.2, 3.5, 3.5, 3.5, 3.6, 3.5, 3.9, 4.6, 5.4, 6.0, 6.5, 7.1, 7.3, 7.3, 7.1, 6.3, 6.2, 6.1, 5.9, 5.8, 6.3, 7.1, 8.1, 8.8, 9.2, 9.1, 9.3, 9.2, 9.3, 8.9, 9.5, 9.8, 10.6, 11.5, 11.9, 12.9, 11.9, 11.7, 10.6, 10.7, 11.2, 9.9, 9.0, 8.9, 8.3, 8.6, 8.5, 8.5, 8.6, 8.8, 8.7, 8.7, 8.8, 9.1, 9.1, 8.8, 9.7, 10.6, 11.7, 9.7, 11.2, 11.1, 9.6, 8.7, 9.0, 8.8, 7.5, 7.3, 7.5, 6.5, 4.3, 4.6, 3.5, 4.3, 3.3, 2.4, 3.5, 4.1, 5.2, 5.6, 5.9, 6.3, 6.8, 7.1, 7.4, 7.5, 7.4, 6.5, 5.9, 5.6, 4.4, 2.9, 2.5, 3.0, 3.2, 2.2, 1.7, 2.3, 2.1, 2.3, 2.7, 3.8, 4.2, 5.9, 6.8, 9.0, 9.4, 10.9, 10.4, 10.2, 7.9, 5.5, 4.7, 2.4, 5.1, 5.1, 4.5, 4.7, 4.0, 4.5, 4.9, 4.2, 4.5, 5.7, 5.0, 5.3, 6.9, 7.9, 9.2, 10.3, 11.6, 12.4, 11.6, 10.8, 9.6, 9.1, 8.8, 9.5, 9.9, 9.9, 9.2, 9.2, 9.1, 9.0, 9.6, 10.2, 10.7, 10.4, 10.3, 10.3, 10.4, 10.7, 11.0, 11.5, 11.4, 11.5, 11.5, 11.5, 11.2, 11.3, 10.9, 10.4, 10.6, 10.2, 9.9, 9.9, 9.5, 9.3, 9.0, 8.9, 8.8, 8.7, 8.5, 8.6, 8.5, 8.9, 8.9, 8.9, 9.0, 8.7, 8.8, 8.7, 8.6, 8.3, 8.5, 8.1, 7.5, 8.0, 8.0, 7.8, 7.6, 7.2, 6.5, 6.4, 6.4, 6.6, 6.6, 6.9, 6.8, 6.8, 7.3, 9.2, 10.5, 10.7, 10.3, 10.2, 8.5, 7.7, 6.4, 5.8, 6.8, 7.2, 7.0, 6.6, 6.7, 5.6, 6.1, 6.2, 5.0, 3.9, 3.4, 3.0, 4.1, 6.4, 8.7, 9.6, 10.8, 10.8, 10.2, 10.3, 7.4, 5.4, 4.4, 2.9, 2.0, 1.2, 1.6, 1.1, 0.9, 1.2, 2.7, 3.3, 4.0, 4.0, 4.8, 5.0, 5.1, 5.1, 5.5, 5.8, 6.7, 7.1, 7.7, 7.8, 7.5, 7.1, 6.6, 4.1, 5.1, 5.6, 5.4, 4.3, 2.8, 3.8, 3.7, 4.1, 4.4, 3.8, 3.8, 3.9, 3.9, 5.5, 6.1, 6.4, 7.2, 7.2, 7.3, 7.1, 6.9, 6.6, 6.1, 5.9, 6.4, 5.0, 4.4, 2.7, 1.4, 3.5, 3.1, 2.0, 2.2, 1.8, 1.0, 1.7, 3.0, 5.1, 7.1, 7.1, 7.8, 7.8, 8.1, 8.2, 8.2, 8.6, 7.9, 7.4, 7.4, 7.3, 7.1, 7.1, 7.0, 7.5, 6.7, 7.0, 6.7, 6.6, 4.8, 4.2, 3.0, 5.1, 6.7, 7.7, 8.0, 8.1, 7.8, 7.4, 6.0, 5.0, 5.0, 4.2, 2.6, 1.4, 0.7, 0.8, 1.6, 1.3, 1.6, 1.6, 0.5, -0.1, 1.4, 1.6, 2.6, 4.7, 5.6, 5.7, 6.3, 7.3, 7.7, 6.1, 6.3, 5.3, 3.4, 3.3, 4.2, 5.8, 6.7, 6.2, 6.4, 7.3, 7.2, 7.9, 7.8, 7.2, 8.1, 5.3, 6.1, 8.1, 11.1, 9.9, 10.3, 10.2, 10.1, 10.0, 9.5, 9.1, 9.6, 8.8, 8.9, 8.8, 8.7, 8.6, 8.6, 8.1, 7.8, 7.6, 7.4, 8.2, 8.2, 9.5, 9.1, 9.0, 9.1, 9.6, 9.7, 9.9, 10.5, 10.4, 9.8, 9.7, 9.4, 9.1, 8.2, 7.6, 7.8, 7.8, 6.1, 6.0, 6.8, 7.2, 7.0, 7.7, 7.8, 7.5, 7.5, 8.2, 8.4, 8.7, 9.3, 9.2, 8.9, 8.6, 8.2, 6.1, 4.9, 4.4, 3.9, 3.5, 3.4, 2.4, 0.8, 0.8, 0.4, 0.3, -0.5, -0.4, -0.3, -0.4, 0.8, 3.0, 3.3, 3.9, 4.6, 5.4, 5.7, 4.2, 2.8, 1.6, 0.8, 1.7, 1.6, 2.1, 3.0, 3.7, 2.8, 4.5, 4.1, 4.6, 5.1, 5.0, 5.1, 5.8, 6.9, 6.9, 7.7, 7.6, 7.3, 7.3, 7.6, 7.8, 7.5, 7.2, 7.3, 7.1, 7.1, 7.0, 6.3, 6.3, 5.5, 6.0, 5.7, 5.6, 5.9, 6.1, 6.0, 6.0, 5.7, 6.1, 7.8, 7.8, 8.3, 8.4, 8.4, 7.4, 6.0, 5.3, 5.0, 4.8, 4.7, 4.8, 4.9, 5.0, 5.0, 4.9, 4.6, 4.5, 4.5, 4.4, 4.3, 4.5, 4.9, 4.9, 5.2, 5.5, 5.6, 5.8, 5.9, 5.7, 5.3, 5.3, 5.0, 4.4, 4.7, 4.8, 3.9, 4.5, 4.3, 4.2, 3.8, 2.3, 1.2, 0.7, 1.8, 2.9, 3.9, 4.8, 5.4, 6.2, 7.0, 7.0, 7.3, 7.6, 7.2, 7.0, 6.4, 6.5, 6.2, 4.3, 4.9, 4.8, 4.7, 5.3, 5.4, 5.7, 6.1, 5.9, 5.7, 5.6, 6.2, 6.3, 7.6, 8.7, 9.9, 10.5, 10.4, 9.3, 8.7, 8.5, 7.9, 8.4, 8.1, 8.4, 7.6, 6.7, 6.1, 5.4, 4.3, 4.0, 3.3, 2.6, 2.2, 2.0, 2.7, 3.9, 5.8, 7.3, 8.6, 10.0, 8.8, 8.0, 5.4, 5.4, 4.7, 3.0, 3.3, 2.7, 3.2, 3.6, 4.3, 4.8, 5.0, 4.1, 3.1, 2.8, 3.1, 2.9, 2.9, 2.8, 3.4, 4.0, 4.4, 4.5, 4.5, 4.9, 4.5, 3.7, 3.4, 2.8, 2.5, 1.1, 0.8, 0.1, 0.0, 1.2, 1.6, 3.2, 3.5, 3.8, 4.0, 4.2, 4.7, 5.0, 5.4, 6.0, 6.4, 6.6, 6.4, 6.2, 5.9, 5.8, 5.8, 5.7, 5.7, 5.5, 5.5, 5.6, 5.5, 5.5, 5.3, 5.2, 5.3, 5.2, 5.0, 5.2, 5.1, 5.2, 5.2, 5.3, 5.4, 5.4, 5.4, 5.5, 5.2, 5.0, 4.9, 4.8, 4.5, 4.3, 4.3, 4.3, 4.2, 4.0, 3.9, 3.9, 3.6, 3.5, 3.1, 2.9, 3.0, 3.4, 3.7, 4.0, 4.3, 4.4, 4.8, 4.8, 5.1, 4.2, 3.4, 2.2, 1.7, 1.3, -0.1, -1.0, -1.6, -1.8, -1.9, -2.3, 0.4, -1.1, -1.1, -1.2, -1.2, 0.8, 2.2, 3.3, 4.0, 3.9, 3.6, 2.8, 1.7, 1.3, 0.2, 0.4, 0.6, 0.3, -1.8, -2.9, -3.7, -4.0, -3.9, -4.5, -5.0, -3.8, -3.5, -4.6, -4.3, -2.1, 0.0, 1.3, 1.8, 3.3, 2.3, 1.8, 0.3, -1.4, -2.7, -3.2, -3.7, -4.0, -3.6, -3.2, -2.7, -2.4, -2.3, -2.8, -2.7, -3.1, -3.8, -3.7, -3.8, -3.5, -2.8, -2.4, -1.7, -1.3, -1.2, -1.6, -2.2, -2.5, -2.5, -2.5, -2.8, -2.6, -3.2, -3.3, -3.5, -3.5, -3.6, -3.9, -3.4, -4.3, -4.2, -4.8, -4.6, -3.2, -2.4, -1.5, -0.6, -0.5, -0.6, -0.7, -2.0, -2.4, -2.8, -3.5, -3.3, -3.6, -3.7, -4.0, -4.4, -5.5, -5.4, -5.2, -5.4, -5.4, -5.3, -5.4, -5.1, -4.4, -3.2, -2.2, -1.5, -0.7, -0.9, -1.7, -2.7, -3.1, -3.5, -3.6, -4.3, -3.9, -5.3, -4.9, -4.9, -6.0, -5.3, -7.3, -5.1, -4.6, -4.4, -4.0, -3.7, -3.1, -2.5, -2.0, -0.3, -0.4, -0.5, -0.8, -1.5, -1.8, -1.8, -2.6, -3.2, -3.4, -3.2, -3.3, -3.1, -3.1, -3.1, -3.0, -2.7, -2.8, -2.4, -3.0, -2.5, -1.6, -0.6, 0.1, 1.7, 1.4, 2.0, 2.2, 1.5, 0.8, 0.6, 0.2, -0.1, 0.1, 0.2, -0.1, 0.0, 0.1, 0.1, 0.0, 0.2, -0.1, -0.3, -0.6, -0.3, 0.3, 2.0, 3.2, 5.2, 4.9, 4.1, 3.4, 1.3, 1.3, 0.4, 0.1, -0.9, -1.2, -1.3, -0.2, 0.2, 0.7, 0.8, 1.0, 1.0, 0.6, 1.3, 1.3, 1.0, 1.8, 2.2, 2.5, 2.7, 2.6, 2.5, 2.4, 2.0, 1.8, 2.0, 1.8, 2.5, 4.6, 4.6, 4.3, 4.6, 4.1, 4.7, 5.8, 5.7, 5.1, 4.8, 5.4, 6.0, 6.3, 6.9, 8.2, 8.4, 8.1, 7.7, 7.2, 7.4, 6.2, 5.9, 6.7, 6.7, 6.4, 5.9, 5.3, 6.0, 6.5, 6.3, 5.8, 6.5, 6.2, 5.4, 5.4, 5.1, 6.3, 6.5, 6.2, 5.4, 5.1, 4.7, 4.5, 4.1, 3.6, 3.2, 3.1, 3.0, 2.8, 2.9, 2.6, 2.2, 2.1, 2.1, 2.0, 2.1, 2.1, 2.1, 2.1, 2.1, 2.2, 2.3, 2.4, 2.6, 2.8, 2.6, 2.3, 2.1, 1.8, 0.8, -0.4, -1.3, -1.6, -1.9, -1.9, -2.7, -2.4, -3.4, -1.7, -1.3, -1.2, -1.1, -2.2, -2.0, 1.6, 2.3, 3.3, 4.2, 5.3, 4.1, 2.3, 0.9, -0.7, -1.4, -2.2, -2.5, -2.4, -3.2, -2.9, -3.0, -3.7, -3.6, -3.4, -2.2, -1.6, -1.1, -0.8, -0.7, 0.4, 2.1, 2.4, 2.2, 2.3, 2.4, 2.4, 2.2, 2.5, 2.6, 3.0, 3.1, 3.3, 3.5, 4.0, 4.0, 4.8, 5.1, 5.2, 5.6, 5.7, 5.9, 5.9, 6.0, 6.3, 6.6, 6.8, 7.2, 7.6, 7.6, 7.3, 7.2, 7.2, 7.3, 7.2, 7.4, 7.5, 7.6, 7.6, 6.8, 6.8, 6.8, 6.6, 6.7, 7.2, 7.2, 7.9, 8.2, 8.4, 8.7, 8.9, 9.2, 9.2, 9.3, 10.2, 10.4, 10.4, 10.9, 11.3, 11.4, 11.8, 12.2, 12.0, 11.8, 11.4, 11.2, 10.7, 10.7, 10.6, 10.3, 9.6, 9.0, 9.1, 9.2, 9.6, 10.0, 10.5, 10.6, 9.7, 9.4, 9.4, 9.0, 8.3, 7.3, 8.1, 7.7, 8.0, 8.0, 7.6, 8.3, 8.5, 8.3, 8.4, 8.9, 8.6, 8.3, 8.8, 9.1, 10.5, 11.4, 11.2, 11.4, 10.9, 10.0, 10.0, 10.1, 9.9, 9.6, 9.9, 9.4, 9.7, 9.5, 9.0, 9.2, 9.0, 8.4, 8.3, 8.2, 7.9, 7.8, 8.0, 8.3, 8.9, 8.8, 9.1, 9.2, 8.9, 8.2, 7.8, 7.4, 7.0, 7.1, 7.5, 7.5, 7.5, 7.4, 7.1, 6.9, 6.7, 6.6, 5.9, 4.9, 6.0, 5.5, 6.7, 7.2, 7.3, 7.3, 7.2, 7.4, 7.9, 8.1, 8.2, 8.4, 8.2, 8.3, 8.4, 6.6, 4.1, 0.8, -1.6, -3.3, -2.8, -2.2, -1.2, -0.5, -0.1, -0.5, -0.3, -0.2, 0.0, 0.1, 0.3, 0.3, 0.2, 0.0, -0.1, -0.1, -0.1, -0.2, -0.3, -0.3, -0.1, 0.0, 0.0, -0.2, -0.1, -0.1, -0.2, -0.3, -0.4, -0.4, -0.4, -0.3, 0.3, 0.5, 0.6, 1.0, 1.6, 1.5, 1.1, 1.4, 1.6, 1.8, 1.8, 1.9, 1.9, 2.0, 1.6, 1.8, 1.8, 2.2, 2.2, 2.1, 0.8, 0.0, 1.4, 3.1, 4.8, 6.2, 6.1, 6.2, 4.6, 3.0, 1.5, 0.5, -0.1, 0.4, 1.6, -0.2, -1.3, -1.9, -2.9, -1.0, -0.7, 1.1, 0.0, -0.5, 0.0, 1.3, 2.3, 3.2, 4.4, 4.9, 5.8, 6.3, 6.1, 6.6, 6.9, 7.6, 7.1, 6.5, 8.0, 7.8, 8.6, 9.5, 12.2, 11.9, 11.1, 10.9, 10.4, 10.3, 9.7, 9.6, 10.2, 10.8, 10.8, 11.1, 11.1, 10.9, 10.4, 9.5, 7.6, 7.2, 8.0, 8.5, 9.2, 8.7, 7.9; 
}